module flop_with_mux(
  input clk,
  input valid,
  input d0,
  input d1,
  input sel,
  output reg q
);

always @(posedge clk) begin
  if (valid) begin
    q <= (sel ? d1 : d0);
  end
end

endmodule

  module ping_buffer (
  input [40-1:0] data_in,
  output [40-1:0] data_out,
  input load_unload, //0 for load (left to right), 1 for unload (top to bottom)
  input valid,
  input clk);

  wire [40-1:0] data_out_internal;
  assign data_out = data_out_internal & {40{load_unload}};
  
wire q_0_0;
wire q_0_1;
wire q_0_2;
wire q_0_3;
wire q_0_4;
wire q_0_5;
wire q_0_6;
wire q_0_7;
wire q_0_8;
wire q_0_9;
wire q_0_10;
wire q_0_11;
wire q_0_12;
wire q_0_13;
wire q_0_14;
wire q_0_15;
wire q_0_16;
wire q_0_17;
wire q_0_18;
wire q_0_19;
wire q_0_20;
wire q_0_21;
wire q_0_22;
wire q_0_23;
wire q_0_24;
wire q_0_25;
wire q_0_26;
wire q_0_27;
wire q_0_28;
wire q_0_29;
wire q_0_30;
wire q_0_31;
wire q_0_32;
wire q_0_33;
wire q_0_34;
wire q_0_35;
wire q_0_36;
wire q_0_37;
wire q_0_38;
wire q_0_39;
wire q_1_0;
wire q_1_1;
wire q_1_2;
wire q_1_3;
wire q_1_4;
wire q_1_5;
wire q_1_6;
wire q_1_7;
wire q_1_8;
wire q_1_9;
wire q_1_10;
wire q_1_11;
wire q_1_12;
wire q_1_13;
wire q_1_14;
wire q_1_15;
wire q_1_16;
wire q_1_17;
wire q_1_18;
wire q_1_19;
wire q_1_20;
wire q_1_21;
wire q_1_22;
wire q_1_23;
wire q_1_24;
wire q_1_25;
wire q_1_26;
wire q_1_27;
wire q_1_28;
wire q_1_29;
wire q_1_30;
wire q_1_31;
wire q_1_32;
wire q_1_33;
wire q_1_34;
wire q_1_35;
wire q_1_36;
wire q_1_37;
wire q_1_38;
wire q_1_39;
wire q_2_0;
wire q_2_1;
wire q_2_2;
wire q_2_3;
wire q_2_4;
wire q_2_5;
wire q_2_6;
wire q_2_7;
wire q_2_8;
wire q_2_9;
wire q_2_10;
wire q_2_11;
wire q_2_12;
wire q_2_13;
wire q_2_14;
wire q_2_15;
wire q_2_16;
wire q_2_17;
wire q_2_18;
wire q_2_19;
wire q_2_20;
wire q_2_21;
wire q_2_22;
wire q_2_23;
wire q_2_24;
wire q_2_25;
wire q_2_26;
wire q_2_27;
wire q_2_28;
wire q_2_29;
wire q_2_30;
wire q_2_31;
wire q_2_32;
wire q_2_33;
wire q_2_34;
wire q_2_35;
wire q_2_36;
wire q_2_37;
wire q_2_38;
wire q_2_39;
wire q_3_0;
wire q_3_1;
wire q_3_2;
wire q_3_3;
wire q_3_4;
wire q_3_5;
wire q_3_6;
wire q_3_7;
wire q_3_8;
wire q_3_9;
wire q_3_10;
wire q_3_11;
wire q_3_12;
wire q_3_13;
wire q_3_14;
wire q_3_15;
wire q_3_16;
wire q_3_17;
wire q_3_18;
wire q_3_19;
wire q_3_20;
wire q_3_21;
wire q_3_22;
wire q_3_23;
wire q_3_24;
wire q_3_25;
wire q_3_26;
wire q_3_27;
wire q_3_28;
wire q_3_29;
wire q_3_30;
wire q_3_31;
wire q_3_32;
wire q_3_33;
wire q_3_34;
wire q_3_35;
wire q_3_36;
wire q_3_37;
wire q_3_38;
wire q_3_39;
wire q_4_0;
wire q_4_1;
wire q_4_2;
wire q_4_3;
wire q_4_4;
wire q_4_5;
wire q_4_6;
wire q_4_7;
wire q_4_8;
wire q_4_9;
wire q_4_10;
wire q_4_11;
wire q_4_12;
wire q_4_13;
wire q_4_14;
wire q_4_15;
wire q_4_16;
wire q_4_17;
wire q_4_18;
wire q_4_19;
wire q_4_20;
wire q_4_21;
wire q_4_22;
wire q_4_23;
wire q_4_24;
wire q_4_25;
wire q_4_26;
wire q_4_27;
wire q_4_28;
wire q_4_29;
wire q_4_30;
wire q_4_31;
wire q_4_32;
wire q_4_33;
wire q_4_34;
wire q_4_35;
wire q_4_36;
wire q_4_37;
wire q_4_38;
wire q_4_39;
wire q_5_0;
wire q_5_1;
wire q_5_2;
wire q_5_3;
wire q_5_4;
wire q_5_5;
wire q_5_6;
wire q_5_7;
wire q_5_8;
wire q_5_9;
wire q_5_10;
wire q_5_11;
wire q_5_12;
wire q_5_13;
wire q_5_14;
wire q_5_15;
wire q_5_16;
wire q_5_17;
wire q_5_18;
wire q_5_19;
wire q_5_20;
wire q_5_21;
wire q_5_22;
wire q_5_23;
wire q_5_24;
wire q_5_25;
wire q_5_26;
wire q_5_27;
wire q_5_28;
wire q_5_29;
wire q_5_30;
wire q_5_31;
wire q_5_32;
wire q_5_33;
wire q_5_34;
wire q_5_35;
wire q_5_36;
wire q_5_37;
wire q_5_38;
wire q_5_39;
wire q_6_0;
wire q_6_1;
wire q_6_2;
wire q_6_3;
wire q_6_4;
wire q_6_5;
wire q_6_6;
wire q_6_7;
wire q_6_8;
wire q_6_9;
wire q_6_10;
wire q_6_11;
wire q_6_12;
wire q_6_13;
wire q_6_14;
wire q_6_15;
wire q_6_16;
wire q_6_17;
wire q_6_18;
wire q_6_19;
wire q_6_20;
wire q_6_21;
wire q_6_22;
wire q_6_23;
wire q_6_24;
wire q_6_25;
wire q_6_26;
wire q_6_27;
wire q_6_28;
wire q_6_29;
wire q_6_30;
wire q_6_31;
wire q_6_32;
wire q_6_33;
wire q_6_34;
wire q_6_35;
wire q_6_36;
wire q_6_37;
wire q_6_38;
wire q_6_39;
wire q_7_0;
wire q_7_1;
wire q_7_2;
wire q_7_3;
wire q_7_4;
wire q_7_5;
wire q_7_6;
wire q_7_7;
wire q_7_8;
wire q_7_9;
wire q_7_10;
wire q_7_11;
wire q_7_12;
wire q_7_13;
wire q_7_14;
wire q_7_15;
wire q_7_16;
wire q_7_17;
wire q_7_18;
wire q_7_19;
wire q_7_20;
wire q_7_21;
wire q_7_22;
wire q_7_23;
wire q_7_24;
wire q_7_25;
wire q_7_26;
wire q_7_27;
wire q_7_28;
wire q_7_29;
wire q_7_30;
wire q_7_31;
wire q_7_32;
wire q_7_33;
wire q_7_34;
wire q_7_35;
wire q_7_36;
wire q_7_37;
wire q_7_38;
wire q_7_39;
wire q_8_0;
wire q_8_1;
wire q_8_2;
wire q_8_3;
wire q_8_4;
wire q_8_5;
wire q_8_6;
wire q_8_7;
wire q_8_8;
wire q_8_9;
wire q_8_10;
wire q_8_11;
wire q_8_12;
wire q_8_13;
wire q_8_14;
wire q_8_15;
wire q_8_16;
wire q_8_17;
wire q_8_18;
wire q_8_19;
wire q_8_20;
wire q_8_21;
wire q_8_22;
wire q_8_23;
wire q_8_24;
wire q_8_25;
wire q_8_26;
wire q_8_27;
wire q_8_28;
wire q_8_29;
wire q_8_30;
wire q_8_31;
wire q_8_32;
wire q_8_33;
wire q_8_34;
wire q_8_35;
wire q_8_36;
wire q_8_37;
wire q_8_38;
wire q_8_39;
wire q_9_0;
wire q_9_1;
wire q_9_2;
wire q_9_3;
wire q_9_4;
wire q_9_5;
wire q_9_6;
wire q_9_7;
wire q_9_8;
wire q_9_9;
wire q_9_10;
wire q_9_11;
wire q_9_12;
wire q_9_13;
wire q_9_14;
wire q_9_15;
wire q_9_16;
wire q_9_17;
wire q_9_18;
wire q_9_19;
wire q_9_20;
wire q_9_21;
wire q_9_22;
wire q_9_23;
wire q_9_24;
wire q_9_25;
wire q_9_26;
wire q_9_27;
wire q_9_28;
wire q_9_29;
wire q_9_30;
wire q_9_31;
wire q_9_32;
wire q_9_33;
wire q_9_34;
wire q_9_35;
wire q_9_36;
wire q_9_37;
wire q_9_38;
wire q_9_39;
wire q_10_0;
wire q_10_1;
wire q_10_2;
wire q_10_3;
wire q_10_4;
wire q_10_5;
wire q_10_6;
wire q_10_7;
wire q_10_8;
wire q_10_9;
wire q_10_10;
wire q_10_11;
wire q_10_12;
wire q_10_13;
wire q_10_14;
wire q_10_15;
wire q_10_16;
wire q_10_17;
wire q_10_18;
wire q_10_19;
wire q_10_20;
wire q_10_21;
wire q_10_22;
wire q_10_23;
wire q_10_24;
wire q_10_25;
wire q_10_26;
wire q_10_27;
wire q_10_28;
wire q_10_29;
wire q_10_30;
wire q_10_31;
wire q_10_32;
wire q_10_33;
wire q_10_34;
wire q_10_35;
wire q_10_36;
wire q_10_37;
wire q_10_38;
wire q_10_39;
wire q_11_0;
wire q_11_1;
wire q_11_2;
wire q_11_3;
wire q_11_4;
wire q_11_5;
wire q_11_6;
wire q_11_7;
wire q_11_8;
wire q_11_9;
wire q_11_10;
wire q_11_11;
wire q_11_12;
wire q_11_13;
wire q_11_14;
wire q_11_15;
wire q_11_16;
wire q_11_17;
wire q_11_18;
wire q_11_19;
wire q_11_20;
wire q_11_21;
wire q_11_22;
wire q_11_23;
wire q_11_24;
wire q_11_25;
wire q_11_26;
wire q_11_27;
wire q_11_28;
wire q_11_29;
wire q_11_30;
wire q_11_31;
wire q_11_32;
wire q_11_33;
wire q_11_34;
wire q_11_35;
wire q_11_36;
wire q_11_37;
wire q_11_38;
wire q_11_39;
wire q_12_0;
wire q_12_1;
wire q_12_2;
wire q_12_3;
wire q_12_4;
wire q_12_5;
wire q_12_6;
wire q_12_7;
wire q_12_8;
wire q_12_9;
wire q_12_10;
wire q_12_11;
wire q_12_12;
wire q_12_13;
wire q_12_14;
wire q_12_15;
wire q_12_16;
wire q_12_17;
wire q_12_18;
wire q_12_19;
wire q_12_20;
wire q_12_21;
wire q_12_22;
wire q_12_23;
wire q_12_24;
wire q_12_25;
wire q_12_26;
wire q_12_27;
wire q_12_28;
wire q_12_29;
wire q_12_30;
wire q_12_31;
wire q_12_32;
wire q_12_33;
wire q_12_34;
wire q_12_35;
wire q_12_36;
wire q_12_37;
wire q_12_38;
wire q_12_39;
wire q_13_0;
wire q_13_1;
wire q_13_2;
wire q_13_3;
wire q_13_4;
wire q_13_5;
wire q_13_6;
wire q_13_7;
wire q_13_8;
wire q_13_9;
wire q_13_10;
wire q_13_11;
wire q_13_12;
wire q_13_13;
wire q_13_14;
wire q_13_15;
wire q_13_16;
wire q_13_17;
wire q_13_18;
wire q_13_19;
wire q_13_20;
wire q_13_21;
wire q_13_22;
wire q_13_23;
wire q_13_24;
wire q_13_25;
wire q_13_26;
wire q_13_27;
wire q_13_28;
wire q_13_29;
wire q_13_30;
wire q_13_31;
wire q_13_32;
wire q_13_33;
wire q_13_34;
wire q_13_35;
wire q_13_36;
wire q_13_37;
wire q_13_38;
wire q_13_39;
wire q_14_0;
wire q_14_1;
wire q_14_2;
wire q_14_3;
wire q_14_4;
wire q_14_5;
wire q_14_6;
wire q_14_7;
wire q_14_8;
wire q_14_9;
wire q_14_10;
wire q_14_11;
wire q_14_12;
wire q_14_13;
wire q_14_14;
wire q_14_15;
wire q_14_16;
wire q_14_17;
wire q_14_18;
wire q_14_19;
wire q_14_20;
wire q_14_21;
wire q_14_22;
wire q_14_23;
wire q_14_24;
wire q_14_25;
wire q_14_26;
wire q_14_27;
wire q_14_28;
wire q_14_29;
wire q_14_30;
wire q_14_31;
wire q_14_32;
wire q_14_33;
wire q_14_34;
wire q_14_35;
wire q_14_36;
wire q_14_37;
wire q_14_38;
wire q_14_39;
wire q_15_0;
wire q_15_1;
wire q_15_2;
wire q_15_3;
wire q_15_4;
wire q_15_5;
wire q_15_6;
wire q_15_7;
wire q_15_8;
wire q_15_9;
wire q_15_10;
wire q_15_11;
wire q_15_12;
wire q_15_13;
wire q_15_14;
wire q_15_15;
wire q_15_16;
wire q_15_17;
wire q_15_18;
wire q_15_19;
wire q_15_20;
wire q_15_21;
wire q_15_22;
wire q_15_23;
wire q_15_24;
wire q_15_25;
wire q_15_26;
wire q_15_27;
wire q_15_28;
wire q_15_29;
wire q_15_30;
wire q_15_31;
wire q_15_32;
wire q_15_33;
wire q_15_34;
wire q_15_35;
wire q_15_36;
wire q_15_37;
wire q_15_38;
wire q_15_39;
wire q_16_0;
wire q_16_1;
wire q_16_2;
wire q_16_3;
wire q_16_4;
wire q_16_5;
wire q_16_6;
wire q_16_7;
wire q_16_8;
wire q_16_9;
wire q_16_10;
wire q_16_11;
wire q_16_12;
wire q_16_13;
wire q_16_14;
wire q_16_15;
wire q_16_16;
wire q_16_17;
wire q_16_18;
wire q_16_19;
wire q_16_20;
wire q_16_21;
wire q_16_22;
wire q_16_23;
wire q_16_24;
wire q_16_25;
wire q_16_26;
wire q_16_27;
wire q_16_28;
wire q_16_29;
wire q_16_30;
wire q_16_31;
wire q_16_32;
wire q_16_33;
wire q_16_34;
wire q_16_35;
wire q_16_36;
wire q_16_37;
wire q_16_38;
wire q_16_39;
wire q_17_0;
wire q_17_1;
wire q_17_2;
wire q_17_3;
wire q_17_4;
wire q_17_5;
wire q_17_6;
wire q_17_7;
wire q_17_8;
wire q_17_9;
wire q_17_10;
wire q_17_11;
wire q_17_12;
wire q_17_13;
wire q_17_14;
wire q_17_15;
wire q_17_16;
wire q_17_17;
wire q_17_18;
wire q_17_19;
wire q_17_20;
wire q_17_21;
wire q_17_22;
wire q_17_23;
wire q_17_24;
wire q_17_25;
wire q_17_26;
wire q_17_27;
wire q_17_28;
wire q_17_29;
wire q_17_30;
wire q_17_31;
wire q_17_32;
wire q_17_33;
wire q_17_34;
wire q_17_35;
wire q_17_36;
wire q_17_37;
wire q_17_38;
wire q_17_39;
wire q_18_0;
wire q_18_1;
wire q_18_2;
wire q_18_3;
wire q_18_4;
wire q_18_5;
wire q_18_6;
wire q_18_7;
wire q_18_8;
wire q_18_9;
wire q_18_10;
wire q_18_11;
wire q_18_12;
wire q_18_13;
wire q_18_14;
wire q_18_15;
wire q_18_16;
wire q_18_17;
wire q_18_18;
wire q_18_19;
wire q_18_20;
wire q_18_21;
wire q_18_22;
wire q_18_23;
wire q_18_24;
wire q_18_25;
wire q_18_26;
wire q_18_27;
wire q_18_28;
wire q_18_29;
wire q_18_30;
wire q_18_31;
wire q_18_32;
wire q_18_33;
wire q_18_34;
wire q_18_35;
wire q_18_36;
wire q_18_37;
wire q_18_38;
wire q_18_39;
wire q_19_0;
wire q_19_1;
wire q_19_2;
wire q_19_3;
wire q_19_4;
wire q_19_5;
wire q_19_6;
wire q_19_7;
wire q_19_8;
wire q_19_9;
wire q_19_10;
wire q_19_11;
wire q_19_12;
wire q_19_13;
wire q_19_14;
wire q_19_15;
wire q_19_16;
wire q_19_17;
wire q_19_18;
wire q_19_19;
wire q_19_20;
wire q_19_21;
wire q_19_22;
wire q_19_23;
wire q_19_24;
wire q_19_25;
wire q_19_26;
wire q_19_27;
wire q_19_28;
wire q_19_29;
wire q_19_30;
wire q_19_31;
wire q_19_32;
wire q_19_33;
wire q_19_34;
wire q_19_35;
wire q_19_36;
wire q_19_37;
wire q_19_38;
wire q_19_39;
wire q_20_0;
wire q_20_1;
wire q_20_2;
wire q_20_3;
wire q_20_4;
wire q_20_5;
wire q_20_6;
wire q_20_7;
wire q_20_8;
wire q_20_9;
wire q_20_10;
wire q_20_11;
wire q_20_12;
wire q_20_13;
wire q_20_14;
wire q_20_15;
wire q_20_16;
wire q_20_17;
wire q_20_18;
wire q_20_19;
wire q_20_20;
wire q_20_21;
wire q_20_22;
wire q_20_23;
wire q_20_24;
wire q_20_25;
wire q_20_26;
wire q_20_27;
wire q_20_28;
wire q_20_29;
wire q_20_30;
wire q_20_31;
wire q_20_32;
wire q_20_33;
wire q_20_34;
wire q_20_35;
wire q_20_36;
wire q_20_37;
wire q_20_38;
wire q_20_39;
wire q_21_0;
wire q_21_1;
wire q_21_2;
wire q_21_3;
wire q_21_4;
wire q_21_5;
wire q_21_6;
wire q_21_7;
wire q_21_8;
wire q_21_9;
wire q_21_10;
wire q_21_11;
wire q_21_12;
wire q_21_13;
wire q_21_14;
wire q_21_15;
wire q_21_16;
wire q_21_17;
wire q_21_18;
wire q_21_19;
wire q_21_20;
wire q_21_21;
wire q_21_22;
wire q_21_23;
wire q_21_24;
wire q_21_25;
wire q_21_26;
wire q_21_27;
wire q_21_28;
wire q_21_29;
wire q_21_30;
wire q_21_31;
wire q_21_32;
wire q_21_33;
wire q_21_34;
wire q_21_35;
wire q_21_36;
wire q_21_37;
wire q_21_38;
wire q_21_39;
wire q_22_0;
wire q_22_1;
wire q_22_2;
wire q_22_3;
wire q_22_4;
wire q_22_5;
wire q_22_6;
wire q_22_7;
wire q_22_8;
wire q_22_9;
wire q_22_10;
wire q_22_11;
wire q_22_12;
wire q_22_13;
wire q_22_14;
wire q_22_15;
wire q_22_16;
wire q_22_17;
wire q_22_18;
wire q_22_19;
wire q_22_20;
wire q_22_21;
wire q_22_22;
wire q_22_23;
wire q_22_24;
wire q_22_25;
wire q_22_26;
wire q_22_27;
wire q_22_28;
wire q_22_29;
wire q_22_30;
wire q_22_31;
wire q_22_32;
wire q_22_33;
wire q_22_34;
wire q_22_35;
wire q_22_36;
wire q_22_37;
wire q_22_38;
wire q_22_39;
wire q_23_0;
wire q_23_1;
wire q_23_2;
wire q_23_3;
wire q_23_4;
wire q_23_5;
wire q_23_6;
wire q_23_7;
wire q_23_8;
wire q_23_9;
wire q_23_10;
wire q_23_11;
wire q_23_12;
wire q_23_13;
wire q_23_14;
wire q_23_15;
wire q_23_16;
wire q_23_17;
wire q_23_18;
wire q_23_19;
wire q_23_20;
wire q_23_21;
wire q_23_22;
wire q_23_23;
wire q_23_24;
wire q_23_25;
wire q_23_26;
wire q_23_27;
wire q_23_28;
wire q_23_29;
wire q_23_30;
wire q_23_31;
wire q_23_32;
wire q_23_33;
wire q_23_34;
wire q_23_35;
wire q_23_36;
wire q_23_37;
wire q_23_38;
wire q_23_39;
wire q_24_0;
wire q_24_1;
wire q_24_2;
wire q_24_3;
wire q_24_4;
wire q_24_5;
wire q_24_6;
wire q_24_7;
wire q_24_8;
wire q_24_9;
wire q_24_10;
wire q_24_11;
wire q_24_12;
wire q_24_13;
wire q_24_14;
wire q_24_15;
wire q_24_16;
wire q_24_17;
wire q_24_18;
wire q_24_19;
wire q_24_20;
wire q_24_21;
wire q_24_22;
wire q_24_23;
wire q_24_24;
wire q_24_25;
wire q_24_26;
wire q_24_27;
wire q_24_28;
wire q_24_29;
wire q_24_30;
wire q_24_31;
wire q_24_32;
wire q_24_33;
wire q_24_34;
wire q_24_35;
wire q_24_36;
wire q_24_37;
wire q_24_38;
wire q_24_39;
wire q_25_0;
wire q_25_1;
wire q_25_2;
wire q_25_3;
wire q_25_4;
wire q_25_5;
wire q_25_6;
wire q_25_7;
wire q_25_8;
wire q_25_9;
wire q_25_10;
wire q_25_11;
wire q_25_12;
wire q_25_13;
wire q_25_14;
wire q_25_15;
wire q_25_16;
wire q_25_17;
wire q_25_18;
wire q_25_19;
wire q_25_20;
wire q_25_21;
wire q_25_22;
wire q_25_23;
wire q_25_24;
wire q_25_25;
wire q_25_26;
wire q_25_27;
wire q_25_28;
wire q_25_29;
wire q_25_30;
wire q_25_31;
wire q_25_32;
wire q_25_33;
wire q_25_34;
wire q_25_35;
wire q_25_36;
wire q_25_37;
wire q_25_38;
wire q_25_39;
wire q_26_0;
wire q_26_1;
wire q_26_2;
wire q_26_3;
wire q_26_4;
wire q_26_5;
wire q_26_6;
wire q_26_7;
wire q_26_8;
wire q_26_9;
wire q_26_10;
wire q_26_11;
wire q_26_12;
wire q_26_13;
wire q_26_14;
wire q_26_15;
wire q_26_16;
wire q_26_17;
wire q_26_18;
wire q_26_19;
wire q_26_20;
wire q_26_21;
wire q_26_22;
wire q_26_23;
wire q_26_24;
wire q_26_25;
wire q_26_26;
wire q_26_27;
wire q_26_28;
wire q_26_29;
wire q_26_30;
wire q_26_31;
wire q_26_32;
wire q_26_33;
wire q_26_34;
wire q_26_35;
wire q_26_36;
wire q_26_37;
wire q_26_38;
wire q_26_39;
wire q_27_0;
wire q_27_1;
wire q_27_2;
wire q_27_3;
wire q_27_4;
wire q_27_5;
wire q_27_6;
wire q_27_7;
wire q_27_8;
wire q_27_9;
wire q_27_10;
wire q_27_11;
wire q_27_12;
wire q_27_13;
wire q_27_14;
wire q_27_15;
wire q_27_16;
wire q_27_17;
wire q_27_18;
wire q_27_19;
wire q_27_20;
wire q_27_21;
wire q_27_22;
wire q_27_23;
wire q_27_24;
wire q_27_25;
wire q_27_26;
wire q_27_27;
wire q_27_28;
wire q_27_29;
wire q_27_30;
wire q_27_31;
wire q_27_32;
wire q_27_33;
wire q_27_34;
wire q_27_35;
wire q_27_36;
wire q_27_37;
wire q_27_38;
wire q_27_39;
wire q_28_0;
wire q_28_1;
wire q_28_2;
wire q_28_3;
wire q_28_4;
wire q_28_5;
wire q_28_6;
wire q_28_7;
wire q_28_8;
wire q_28_9;
wire q_28_10;
wire q_28_11;
wire q_28_12;
wire q_28_13;
wire q_28_14;
wire q_28_15;
wire q_28_16;
wire q_28_17;
wire q_28_18;
wire q_28_19;
wire q_28_20;
wire q_28_21;
wire q_28_22;
wire q_28_23;
wire q_28_24;
wire q_28_25;
wire q_28_26;
wire q_28_27;
wire q_28_28;
wire q_28_29;
wire q_28_30;
wire q_28_31;
wire q_28_32;
wire q_28_33;
wire q_28_34;
wire q_28_35;
wire q_28_36;
wire q_28_37;
wire q_28_38;
wire q_28_39;
wire q_29_0;
wire q_29_1;
wire q_29_2;
wire q_29_3;
wire q_29_4;
wire q_29_5;
wire q_29_6;
wire q_29_7;
wire q_29_8;
wire q_29_9;
wire q_29_10;
wire q_29_11;
wire q_29_12;
wire q_29_13;
wire q_29_14;
wire q_29_15;
wire q_29_16;
wire q_29_17;
wire q_29_18;
wire q_29_19;
wire q_29_20;
wire q_29_21;
wire q_29_22;
wire q_29_23;
wire q_29_24;
wire q_29_25;
wire q_29_26;
wire q_29_27;
wire q_29_28;
wire q_29_29;
wire q_29_30;
wire q_29_31;
wire q_29_32;
wire q_29_33;
wire q_29_34;
wire q_29_35;
wire q_29_36;
wire q_29_37;
wire q_29_38;
wire q_29_39;
wire q_30_0;
wire q_30_1;
wire q_30_2;
wire q_30_3;
wire q_30_4;
wire q_30_5;
wire q_30_6;
wire q_30_7;
wire q_30_8;
wire q_30_9;
wire q_30_10;
wire q_30_11;
wire q_30_12;
wire q_30_13;
wire q_30_14;
wire q_30_15;
wire q_30_16;
wire q_30_17;
wire q_30_18;
wire q_30_19;
wire q_30_20;
wire q_30_21;
wire q_30_22;
wire q_30_23;
wire q_30_24;
wire q_30_25;
wire q_30_26;
wire q_30_27;
wire q_30_28;
wire q_30_29;
wire q_30_30;
wire q_30_31;
wire q_30_32;
wire q_30_33;
wire q_30_34;
wire q_30_35;
wire q_30_36;
wire q_30_37;
wire q_30_38;
wire q_30_39;
wire q_31_0;
wire q_31_1;
wire q_31_2;
wire q_31_3;
wire q_31_4;
wire q_31_5;
wire q_31_6;
wire q_31_7;
wire q_31_8;
wire q_31_9;
wire q_31_10;
wire q_31_11;
wire q_31_12;
wire q_31_13;
wire q_31_14;
wire q_31_15;
wire q_31_16;
wire q_31_17;
wire q_31_18;
wire q_31_19;
wire q_31_20;
wire q_31_21;
wire q_31_22;
wire q_31_23;
wire q_31_24;
wire q_31_25;
wire q_31_26;
wire q_31_27;
wire q_31_28;
wire q_31_29;
wire q_31_30;
wire q_31_31;
wire q_31_32;
wire q_31_33;
wire q_31_34;
wire q_31_35;
wire q_31_36;
wire q_31_37;
wire q_31_38;
wire q_31_39;
wire q_32_0;
wire q_32_1;
wire q_32_2;
wire q_32_3;
wire q_32_4;
wire q_32_5;
wire q_32_6;
wire q_32_7;
wire q_32_8;
wire q_32_9;
wire q_32_10;
wire q_32_11;
wire q_32_12;
wire q_32_13;
wire q_32_14;
wire q_32_15;
wire q_32_16;
wire q_32_17;
wire q_32_18;
wire q_32_19;
wire q_32_20;
wire q_32_21;
wire q_32_22;
wire q_32_23;
wire q_32_24;
wire q_32_25;
wire q_32_26;
wire q_32_27;
wire q_32_28;
wire q_32_29;
wire q_32_30;
wire q_32_31;
wire q_32_32;
wire q_32_33;
wire q_32_34;
wire q_32_35;
wire q_32_36;
wire q_32_37;
wire q_32_38;
wire q_32_39;
wire q_33_0;
wire q_33_1;
wire q_33_2;
wire q_33_3;
wire q_33_4;
wire q_33_5;
wire q_33_6;
wire q_33_7;
wire q_33_8;
wire q_33_9;
wire q_33_10;
wire q_33_11;
wire q_33_12;
wire q_33_13;
wire q_33_14;
wire q_33_15;
wire q_33_16;
wire q_33_17;
wire q_33_18;
wire q_33_19;
wire q_33_20;
wire q_33_21;
wire q_33_22;
wire q_33_23;
wire q_33_24;
wire q_33_25;
wire q_33_26;
wire q_33_27;
wire q_33_28;
wire q_33_29;
wire q_33_30;
wire q_33_31;
wire q_33_32;
wire q_33_33;
wire q_33_34;
wire q_33_35;
wire q_33_36;
wire q_33_37;
wire q_33_38;
wire q_33_39;
wire q_34_0;
wire q_34_1;
wire q_34_2;
wire q_34_3;
wire q_34_4;
wire q_34_5;
wire q_34_6;
wire q_34_7;
wire q_34_8;
wire q_34_9;
wire q_34_10;
wire q_34_11;
wire q_34_12;
wire q_34_13;
wire q_34_14;
wire q_34_15;
wire q_34_16;
wire q_34_17;
wire q_34_18;
wire q_34_19;
wire q_34_20;
wire q_34_21;
wire q_34_22;
wire q_34_23;
wire q_34_24;
wire q_34_25;
wire q_34_26;
wire q_34_27;
wire q_34_28;
wire q_34_29;
wire q_34_30;
wire q_34_31;
wire q_34_32;
wire q_34_33;
wire q_34_34;
wire q_34_35;
wire q_34_36;
wire q_34_37;
wire q_34_38;
wire q_34_39;
wire q_35_0;
wire q_35_1;
wire q_35_2;
wire q_35_3;
wire q_35_4;
wire q_35_5;
wire q_35_6;
wire q_35_7;
wire q_35_8;
wire q_35_9;
wire q_35_10;
wire q_35_11;
wire q_35_12;
wire q_35_13;
wire q_35_14;
wire q_35_15;
wire q_35_16;
wire q_35_17;
wire q_35_18;
wire q_35_19;
wire q_35_20;
wire q_35_21;
wire q_35_22;
wire q_35_23;
wire q_35_24;
wire q_35_25;
wire q_35_26;
wire q_35_27;
wire q_35_28;
wire q_35_29;
wire q_35_30;
wire q_35_31;
wire q_35_32;
wire q_35_33;
wire q_35_34;
wire q_35_35;
wire q_35_36;
wire q_35_37;
wire q_35_38;
wire q_35_39;
wire q_36_0;
wire q_36_1;
wire q_36_2;
wire q_36_3;
wire q_36_4;
wire q_36_5;
wire q_36_6;
wire q_36_7;
wire q_36_8;
wire q_36_9;
wire q_36_10;
wire q_36_11;
wire q_36_12;
wire q_36_13;
wire q_36_14;
wire q_36_15;
wire q_36_16;
wire q_36_17;
wire q_36_18;
wire q_36_19;
wire q_36_20;
wire q_36_21;
wire q_36_22;
wire q_36_23;
wire q_36_24;
wire q_36_25;
wire q_36_26;
wire q_36_27;
wire q_36_28;
wire q_36_29;
wire q_36_30;
wire q_36_31;
wire q_36_32;
wire q_36_33;
wire q_36_34;
wire q_36_35;
wire q_36_36;
wire q_36_37;
wire q_36_38;
wire q_36_39;
wire q_37_0;
wire q_37_1;
wire q_37_2;
wire q_37_3;
wire q_37_4;
wire q_37_5;
wire q_37_6;
wire q_37_7;
wire q_37_8;
wire q_37_9;
wire q_37_10;
wire q_37_11;
wire q_37_12;
wire q_37_13;
wire q_37_14;
wire q_37_15;
wire q_37_16;
wire q_37_17;
wire q_37_18;
wire q_37_19;
wire q_37_20;
wire q_37_21;
wire q_37_22;
wire q_37_23;
wire q_37_24;
wire q_37_25;
wire q_37_26;
wire q_37_27;
wire q_37_28;
wire q_37_29;
wire q_37_30;
wire q_37_31;
wire q_37_32;
wire q_37_33;
wire q_37_34;
wire q_37_35;
wire q_37_36;
wire q_37_37;
wire q_37_38;
wire q_37_39;
wire q_38_0;
wire q_38_1;
wire q_38_2;
wire q_38_3;
wire q_38_4;
wire q_38_5;
wire q_38_6;
wire q_38_7;
wire q_38_8;
wire q_38_9;
wire q_38_10;
wire q_38_11;
wire q_38_12;
wire q_38_13;
wire q_38_14;
wire q_38_15;
wire q_38_16;
wire q_38_17;
wire q_38_18;
wire q_38_19;
wire q_38_20;
wire q_38_21;
wire q_38_22;
wire q_38_23;
wire q_38_24;
wire q_38_25;
wire q_38_26;
wire q_38_27;
wire q_38_28;
wire q_38_29;
wire q_38_30;
wire q_38_31;
wire q_38_32;
wire q_38_33;
wire q_38_34;
wire q_38_35;
wire q_38_36;
wire q_38_37;
wire q_38_38;
wire q_38_39;
wire q_39_0;
wire q_39_1;
wire q_39_2;
wire q_39_3;
wire q_39_4;
wire q_39_5;
wire q_39_6;
wire q_39_7;
wire q_39_8;
wire q_39_9;
wire q_39_10;
wire q_39_11;
wire q_39_12;
wire q_39_13;
wire q_39_14;
wire q_39_15;
wire q_39_16;
wire q_39_17;
wire q_39_18;
wire q_39_19;
wire q_39_20;
wire q_39_21;
wire q_39_22;
wire q_39_23;
wire q_39_24;
wire q_39_25;
wire q_39_26;
wire q_39_27;
wire q_39_28;
wire q_39_29;
wire q_39_30;
wire q_39_31;
wire q_39_32;
wire q_39_33;
wire q_39_34;
wire q_39_35;
wire q_39_36;
wire q_39_37;
wire q_39_38;
wire q_39_39;

  wire q_0_minus1;
  assign q_0_minus1 = data_in[0];
  

  wire q_1_minus1;
  assign q_1_minus1 = data_in[1];
  

  wire q_2_minus1;
  assign q_2_minus1 = data_in[2];
  

  wire q_3_minus1;
  assign q_3_minus1 = data_in[3];
  

  wire q_4_minus1;
  assign q_4_minus1 = data_in[4];
  

  wire q_5_minus1;
  assign q_5_minus1 = data_in[5];
  

  wire q_6_minus1;
  assign q_6_minus1 = data_in[6];
  

  wire q_7_minus1;
  assign q_7_minus1 = data_in[7];
  

  wire q_8_minus1;
  assign q_8_minus1 = data_in[8];
  

  wire q_9_minus1;
  assign q_9_minus1 = data_in[9];
  

  wire q_10_minus1;
  assign q_10_minus1 = data_in[10];
  

  wire q_11_minus1;
  assign q_11_minus1 = data_in[11];
  

  wire q_12_minus1;
  assign q_12_minus1 = data_in[12];
  

  wire q_13_minus1;
  assign q_13_minus1 = data_in[13];
  

  wire q_14_minus1;
  assign q_14_minus1 = data_in[14];
  

  wire q_15_minus1;
  assign q_15_minus1 = data_in[15];
  

  wire q_16_minus1;
  assign q_16_minus1 = data_in[16];
  

  wire q_17_minus1;
  assign q_17_minus1 = data_in[17];
  

  wire q_18_minus1;
  assign q_18_minus1 = data_in[18];
  

  wire q_19_minus1;
  assign q_19_minus1 = data_in[19];
  

  wire q_20_minus1;
  assign q_20_minus1 = data_in[20];
  

  wire q_21_minus1;
  assign q_21_minus1 = data_in[21];
  

  wire q_22_minus1;
  assign q_22_minus1 = data_in[22];
  

  wire q_23_minus1;
  assign q_23_minus1 = data_in[23];
  

  wire q_24_minus1;
  assign q_24_minus1 = data_in[24];
  

  wire q_25_minus1;
  assign q_25_minus1 = data_in[25];
  

  wire q_26_minus1;
  assign q_26_minus1 = data_in[26];
  

  wire q_27_minus1;
  assign q_27_minus1 = data_in[27];
  

  wire q_28_minus1;
  assign q_28_minus1 = data_in[28];
  

  wire q_29_minus1;
  assign q_29_minus1 = data_in[29];
  

  wire q_30_minus1;
  assign q_30_minus1 = data_in[30];
  

  wire q_31_minus1;
  assign q_31_minus1 = data_in[31];
  

  wire q_32_minus1;
  assign q_32_minus1 = data_in[32];
  

  wire q_33_minus1;
  assign q_33_minus1 = data_in[33];
  

  wire q_34_minus1;
  assign q_34_minus1 = data_in[34];
  

  wire q_35_minus1;
  assign q_35_minus1 = data_in[35];
  

  wire q_36_minus1;
  assign q_36_minus1 = data_in[36];
  

  wire q_37_minus1;
  assign q_37_minus1 = data_in[37];
  

  wire q_38_minus1;
  assign q_38_minus1 = data_in[38];
  

  wire q_39_minus1;
  assign q_39_minus1 = data_in[39];
  

  assign data_out_internal[0] = q_39_0;
  

  assign data_out_internal[1] = q_39_1;
  

  assign data_out_internal[2] = q_39_2;
  

  assign data_out_internal[3] = q_39_3;
  

  assign data_out_internal[4] = q_39_4;
  

  assign data_out_internal[5] = q_39_5;
  

  assign data_out_internal[6] = q_39_6;
  

  assign data_out_internal[7] = q_39_7;
  

  assign data_out_internal[8] = q_39_8;
  

  assign data_out_internal[9] = q_39_9;
  

  assign data_out_internal[10] = q_39_10;
  

  assign data_out_internal[11] = q_39_11;
  

  assign data_out_internal[12] = q_39_12;
  

  assign data_out_internal[13] = q_39_13;
  

  assign data_out_internal[14] = q_39_14;
  

  assign data_out_internal[15] = q_39_15;
  

  assign data_out_internal[16] = q_39_16;
  

  assign data_out_internal[17] = q_39_17;
  

  assign data_out_internal[18] = q_39_18;
  

  assign data_out_internal[19] = q_39_19;
  

  assign data_out_internal[20] = q_39_20;
  

  assign data_out_internal[21] = q_39_21;
  

  assign data_out_internal[22] = q_39_22;
  

  assign data_out_internal[23] = q_39_23;
  

  assign data_out_internal[24] = q_39_24;
  

  assign data_out_internal[25] = q_39_25;
  

  assign data_out_internal[26] = q_39_26;
  

  assign data_out_internal[27] = q_39_27;
  

  assign data_out_internal[28] = q_39_28;
  

  assign data_out_internal[29] = q_39_29;
  

  assign data_out_internal[30] = q_39_30;
  

  assign data_out_internal[31] = q_39_31;
  

  assign data_out_internal[32] = q_39_32;
  

  assign data_out_internal[33] = q_39_33;
  

  assign data_out_internal[34] = q_39_34;
  

  assign data_out_internal[35] = q_39_35;
  

  assign data_out_internal[36] = q_39_36;
  

  assign data_out_internal[37] = q_39_37;
  

  assign data_out_internal[38] = q_39_38;
  

  assign data_out_internal[39] = q_39_39;
  

  wire q_minus1_0;
  assign q_minus1_0 = 1'b0;
  

  wire q_minus1_1;
  assign q_minus1_1 = 1'b0;
  

  wire q_minus1_2;
  assign q_minus1_2 = 1'b0;
  

  wire q_minus1_3;
  assign q_minus1_3 = 1'b0;
  

  wire q_minus1_4;
  assign q_minus1_4 = 1'b0;
  

  wire q_minus1_5;
  assign q_minus1_5 = 1'b0;
  

  wire q_minus1_6;
  assign q_minus1_6 = 1'b0;
  

  wire q_minus1_7;
  assign q_minus1_7 = 1'b0;
  

  wire q_minus1_8;
  assign q_minus1_8 = 1'b0;
  

  wire q_minus1_9;
  assign q_minus1_9 = 1'b0;
  

  wire q_minus1_10;
  assign q_minus1_10 = 1'b0;
  

  wire q_minus1_11;
  assign q_minus1_11 = 1'b0;
  

  wire q_minus1_12;
  assign q_minus1_12 = 1'b0;
  

  wire q_minus1_13;
  assign q_minus1_13 = 1'b0;
  

  wire q_minus1_14;
  assign q_minus1_14 = 1'b0;
  

  wire q_minus1_15;
  assign q_minus1_15 = 1'b0;
  

  wire q_minus1_16;
  assign q_minus1_16 = 1'b0;
  

  wire q_minus1_17;
  assign q_minus1_17 = 1'b0;
  

  wire q_minus1_18;
  assign q_minus1_18 = 1'b0;
  

  wire q_minus1_19;
  assign q_minus1_19 = 1'b0;
  

  wire q_minus1_20;
  assign q_minus1_20 = 1'b0;
  

  wire q_minus1_21;
  assign q_minus1_21 = 1'b0;
  

  wire q_minus1_22;
  assign q_minus1_22 = 1'b0;
  

  wire q_minus1_23;
  assign q_minus1_23 = 1'b0;
  

  wire q_minus1_24;
  assign q_minus1_24 = 1'b0;
  

  wire q_minus1_25;
  assign q_minus1_25 = 1'b0;
  

  wire q_minus1_26;
  assign q_minus1_26 = 1'b0;
  

  wire q_minus1_27;
  assign q_minus1_27 = 1'b0;
  

  wire q_minus1_28;
  assign q_minus1_28 = 1'b0;
  

  wire q_minus1_29;
  assign q_minus1_29 = 1'b0;
  

  wire q_minus1_30;
  assign q_minus1_30 = 1'b0;
  

  wire q_minus1_31;
  assign q_minus1_31 = 1'b0;
  

  wire q_minus1_32;
  assign q_minus1_32 = 1'b0;
  

  wire q_minus1_33;
  assign q_minus1_33 = 1'b0;
  

  wire q_minus1_34;
  assign q_minus1_34 = 1'b0;
  

  wire q_minus1_35;
  assign q_minus1_35 = 1'b0;
  

  wire q_minus1_36;
  assign q_minus1_36 = 1'b0;
  

  wire q_minus1_37;
  assign q_minus1_37 = 1'b0;
  

  wire q_minus1_38;
  assign q_minus1_38 = 1'b0;
  

  wire q_minus1_39;
  assign q_minus1_39 = 1'b0;
  

  flop_with_mux u_0_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_minus1),
    .d1(q_minus1_0),
    .q(q_0_0)
  );
  

  flop_with_mux u_0_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_0),
    .d1(q_minus1_1),
    .q(q_0_1)
  );
  

  flop_with_mux u_0_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_1),
    .d1(q_minus1_2),
    .q(q_0_2)
  );
  

  flop_with_mux u_0_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_2),
    .d1(q_minus1_3),
    .q(q_0_3)
  );
  

  flop_with_mux u_0_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_3),
    .d1(q_minus1_4),
    .q(q_0_4)
  );
  

  flop_with_mux u_0_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_4),
    .d1(q_minus1_5),
    .q(q_0_5)
  );
  

  flop_with_mux u_0_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_5),
    .d1(q_minus1_6),
    .q(q_0_6)
  );
  

  flop_with_mux u_0_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_6),
    .d1(q_minus1_7),
    .q(q_0_7)
  );
  

  flop_with_mux u_0_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_7),
    .d1(q_minus1_8),
    .q(q_0_8)
  );
  

  flop_with_mux u_0_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_8),
    .d1(q_minus1_9),
    .q(q_0_9)
  );
  

  flop_with_mux u_0_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_9),
    .d1(q_minus1_10),
    .q(q_0_10)
  );
  

  flop_with_mux u_0_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_10),
    .d1(q_minus1_11),
    .q(q_0_11)
  );
  

  flop_with_mux u_0_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_11),
    .d1(q_minus1_12),
    .q(q_0_12)
  );
  

  flop_with_mux u_0_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_12),
    .d1(q_minus1_13),
    .q(q_0_13)
  );
  

  flop_with_mux u_0_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_13),
    .d1(q_minus1_14),
    .q(q_0_14)
  );
  

  flop_with_mux u_0_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_14),
    .d1(q_minus1_15),
    .q(q_0_15)
  );
  

  flop_with_mux u_0_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_15),
    .d1(q_minus1_16),
    .q(q_0_16)
  );
  

  flop_with_mux u_0_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_16),
    .d1(q_minus1_17),
    .q(q_0_17)
  );
  

  flop_with_mux u_0_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_17),
    .d1(q_minus1_18),
    .q(q_0_18)
  );
  

  flop_with_mux u_0_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_18),
    .d1(q_minus1_19),
    .q(q_0_19)
  );
  

  flop_with_mux u_0_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_19),
    .d1(q_minus1_20),
    .q(q_0_20)
  );
  

  flop_with_mux u_0_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_20),
    .d1(q_minus1_21),
    .q(q_0_21)
  );
  

  flop_with_mux u_0_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_21),
    .d1(q_minus1_22),
    .q(q_0_22)
  );
  

  flop_with_mux u_0_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_22),
    .d1(q_minus1_23),
    .q(q_0_23)
  );
  

  flop_with_mux u_0_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_23),
    .d1(q_minus1_24),
    .q(q_0_24)
  );
  

  flop_with_mux u_0_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_24),
    .d1(q_minus1_25),
    .q(q_0_25)
  );
  

  flop_with_mux u_0_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_25),
    .d1(q_minus1_26),
    .q(q_0_26)
  );
  

  flop_with_mux u_0_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_26),
    .d1(q_minus1_27),
    .q(q_0_27)
  );
  

  flop_with_mux u_0_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_27),
    .d1(q_minus1_28),
    .q(q_0_28)
  );
  

  flop_with_mux u_0_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_28),
    .d1(q_minus1_29),
    .q(q_0_29)
  );
  

  flop_with_mux u_0_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_29),
    .d1(q_minus1_30),
    .q(q_0_30)
  );
  

  flop_with_mux u_0_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_30),
    .d1(q_minus1_31),
    .q(q_0_31)
  );
  

  flop_with_mux u_0_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_31),
    .d1(q_minus1_32),
    .q(q_0_32)
  );
  

  flop_with_mux u_0_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_32),
    .d1(q_minus1_33),
    .q(q_0_33)
  );
  

  flop_with_mux u_0_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_33),
    .d1(q_minus1_34),
    .q(q_0_34)
  );
  

  flop_with_mux u_0_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_34),
    .d1(q_minus1_35),
    .q(q_0_35)
  );
  

  flop_with_mux u_0_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_35),
    .d1(q_minus1_36),
    .q(q_0_36)
  );
  

  flop_with_mux u_0_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_36),
    .d1(q_minus1_37),
    .q(q_0_37)
  );
  

  flop_with_mux u_0_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_37),
    .d1(q_minus1_38),
    .q(q_0_38)
  );
  

  flop_with_mux u_0_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_38),
    .d1(q_minus1_39),
    .q(q_0_39)
  );
  

  flop_with_mux u_1_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_minus1),
    .d1(q_0_0),
    .q(q_1_0)
  );
  

  flop_with_mux u_1_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_0),
    .d1(q_0_1),
    .q(q_1_1)
  );
  

  flop_with_mux u_1_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_1),
    .d1(q_0_2),
    .q(q_1_2)
  );
  

  flop_with_mux u_1_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_2),
    .d1(q_0_3),
    .q(q_1_3)
  );
  

  flop_with_mux u_1_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_3),
    .d1(q_0_4),
    .q(q_1_4)
  );
  

  flop_with_mux u_1_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_4),
    .d1(q_0_5),
    .q(q_1_5)
  );
  

  flop_with_mux u_1_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_5),
    .d1(q_0_6),
    .q(q_1_6)
  );
  

  flop_with_mux u_1_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_6),
    .d1(q_0_7),
    .q(q_1_7)
  );
  

  flop_with_mux u_1_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_7),
    .d1(q_0_8),
    .q(q_1_8)
  );
  

  flop_with_mux u_1_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_8),
    .d1(q_0_9),
    .q(q_1_9)
  );
  

  flop_with_mux u_1_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_9),
    .d1(q_0_10),
    .q(q_1_10)
  );
  

  flop_with_mux u_1_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_10),
    .d1(q_0_11),
    .q(q_1_11)
  );
  

  flop_with_mux u_1_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_11),
    .d1(q_0_12),
    .q(q_1_12)
  );
  

  flop_with_mux u_1_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_12),
    .d1(q_0_13),
    .q(q_1_13)
  );
  

  flop_with_mux u_1_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_13),
    .d1(q_0_14),
    .q(q_1_14)
  );
  

  flop_with_mux u_1_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_14),
    .d1(q_0_15),
    .q(q_1_15)
  );
  

  flop_with_mux u_1_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_15),
    .d1(q_0_16),
    .q(q_1_16)
  );
  

  flop_with_mux u_1_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_16),
    .d1(q_0_17),
    .q(q_1_17)
  );
  

  flop_with_mux u_1_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_17),
    .d1(q_0_18),
    .q(q_1_18)
  );
  

  flop_with_mux u_1_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_18),
    .d1(q_0_19),
    .q(q_1_19)
  );
  

  flop_with_mux u_1_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_19),
    .d1(q_0_20),
    .q(q_1_20)
  );
  

  flop_with_mux u_1_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_20),
    .d1(q_0_21),
    .q(q_1_21)
  );
  

  flop_with_mux u_1_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_21),
    .d1(q_0_22),
    .q(q_1_22)
  );
  

  flop_with_mux u_1_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_22),
    .d1(q_0_23),
    .q(q_1_23)
  );
  

  flop_with_mux u_1_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_23),
    .d1(q_0_24),
    .q(q_1_24)
  );
  

  flop_with_mux u_1_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_24),
    .d1(q_0_25),
    .q(q_1_25)
  );
  

  flop_with_mux u_1_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_25),
    .d1(q_0_26),
    .q(q_1_26)
  );
  

  flop_with_mux u_1_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_26),
    .d1(q_0_27),
    .q(q_1_27)
  );
  

  flop_with_mux u_1_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_27),
    .d1(q_0_28),
    .q(q_1_28)
  );
  

  flop_with_mux u_1_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_28),
    .d1(q_0_29),
    .q(q_1_29)
  );
  

  flop_with_mux u_1_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_29),
    .d1(q_0_30),
    .q(q_1_30)
  );
  

  flop_with_mux u_1_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_30),
    .d1(q_0_31),
    .q(q_1_31)
  );
  

  flop_with_mux u_1_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_31),
    .d1(q_0_32),
    .q(q_1_32)
  );
  

  flop_with_mux u_1_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_32),
    .d1(q_0_33),
    .q(q_1_33)
  );
  

  flop_with_mux u_1_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_33),
    .d1(q_0_34),
    .q(q_1_34)
  );
  

  flop_with_mux u_1_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_34),
    .d1(q_0_35),
    .q(q_1_35)
  );
  

  flop_with_mux u_1_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_35),
    .d1(q_0_36),
    .q(q_1_36)
  );
  

  flop_with_mux u_1_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_36),
    .d1(q_0_37),
    .q(q_1_37)
  );
  

  flop_with_mux u_1_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_37),
    .d1(q_0_38),
    .q(q_1_38)
  );
  

  flop_with_mux u_1_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_38),
    .d1(q_0_39),
    .q(q_1_39)
  );
  

  flop_with_mux u_2_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_minus1),
    .d1(q_1_0),
    .q(q_2_0)
  );
  

  flop_with_mux u_2_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_0),
    .d1(q_1_1),
    .q(q_2_1)
  );
  

  flop_with_mux u_2_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_1),
    .d1(q_1_2),
    .q(q_2_2)
  );
  

  flop_with_mux u_2_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_2),
    .d1(q_1_3),
    .q(q_2_3)
  );
  

  flop_with_mux u_2_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_3),
    .d1(q_1_4),
    .q(q_2_4)
  );
  

  flop_with_mux u_2_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_4),
    .d1(q_1_5),
    .q(q_2_5)
  );
  

  flop_with_mux u_2_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_5),
    .d1(q_1_6),
    .q(q_2_6)
  );
  

  flop_with_mux u_2_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_6),
    .d1(q_1_7),
    .q(q_2_7)
  );
  

  flop_with_mux u_2_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_7),
    .d1(q_1_8),
    .q(q_2_8)
  );
  

  flop_with_mux u_2_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_8),
    .d1(q_1_9),
    .q(q_2_9)
  );
  

  flop_with_mux u_2_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_9),
    .d1(q_1_10),
    .q(q_2_10)
  );
  

  flop_with_mux u_2_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_10),
    .d1(q_1_11),
    .q(q_2_11)
  );
  

  flop_with_mux u_2_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_11),
    .d1(q_1_12),
    .q(q_2_12)
  );
  

  flop_with_mux u_2_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_12),
    .d1(q_1_13),
    .q(q_2_13)
  );
  

  flop_with_mux u_2_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_13),
    .d1(q_1_14),
    .q(q_2_14)
  );
  

  flop_with_mux u_2_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_14),
    .d1(q_1_15),
    .q(q_2_15)
  );
  

  flop_with_mux u_2_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_15),
    .d1(q_1_16),
    .q(q_2_16)
  );
  

  flop_with_mux u_2_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_16),
    .d1(q_1_17),
    .q(q_2_17)
  );
  

  flop_with_mux u_2_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_17),
    .d1(q_1_18),
    .q(q_2_18)
  );
  

  flop_with_mux u_2_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_18),
    .d1(q_1_19),
    .q(q_2_19)
  );
  

  flop_with_mux u_2_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_19),
    .d1(q_1_20),
    .q(q_2_20)
  );
  

  flop_with_mux u_2_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_20),
    .d1(q_1_21),
    .q(q_2_21)
  );
  

  flop_with_mux u_2_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_21),
    .d1(q_1_22),
    .q(q_2_22)
  );
  

  flop_with_mux u_2_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_22),
    .d1(q_1_23),
    .q(q_2_23)
  );
  

  flop_with_mux u_2_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_23),
    .d1(q_1_24),
    .q(q_2_24)
  );
  

  flop_with_mux u_2_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_24),
    .d1(q_1_25),
    .q(q_2_25)
  );
  

  flop_with_mux u_2_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_25),
    .d1(q_1_26),
    .q(q_2_26)
  );
  

  flop_with_mux u_2_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_26),
    .d1(q_1_27),
    .q(q_2_27)
  );
  

  flop_with_mux u_2_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_27),
    .d1(q_1_28),
    .q(q_2_28)
  );
  

  flop_with_mux u_2_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_28),
    .d1(q_1_29),
    .q(q_2_29)
  );
  

  flop_with_mux u_2_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_29),
    .d1(q_1_30),
    .q(q_2_30)
  );
  

  flop_with_mux u_2_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_30),
    .d1(q_1_31),
    .q(q_2_31)
  );
  

  flop_with_mux u_2_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_31),
    .d1(q_1_32),
    .q(q_2_32)
  );
  

  flop_with_mux u_2_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_32),
    .d1(q_1_33),
    .q(q_2_33)
  );
  

  flop_with_mux u_2_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_33),
    .d1(q_1_34),
    .q(q_2_34)
  );
  

  flop_with_mux u_2_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_34),
    .d1(q_1_35),
    .q(q_2_35)
  );
  

  flop_with_mux u_2_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_35),
    .d1(q_1_36),
    .q(q_2_36)
  );
  

  flop_with_mux u_2_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_36),
    .d1(q_1_37),
    .q(q_2_37)
  );
  

  flop_with_mux u_2_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_37),
    .d1(q_1_38),
    .q(q_2_38)
  );
  

  flop_with_mux u_2_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_38),
    .d1(q_1_39),
    .q(q_2_39)
  );
  

  flop_with_mux u_3_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_minus1),
    .d1(q_2_0),
    .q(q_3_0)
  );
  

  flop_with_mux u_3_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_0),
    .d1(q_2_1),
    .q(q_3_1)
  );
  

  flop_with_mux u_3_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_1),
    .d1(q_2_2),
    .q(q_3_2)
  );
  

  flop_with_mux u_3_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_2),
    .d1(q_2_3),
    .q(q_3_3)
  );
  

  flop_with_mux u_3_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_3),
    .d1(q_2_4),
    .q(q_3_4)
  );
  

  flop_with_mux u_3_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_4),
    .d1(q_2_5),
    .q(q_3_5)
  );
  

  flop_with_mux u_3_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_5),
    .d1(q_2_6),
    .q(q_3_6)
  );
  

  flop_with_mux u_3_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_6),
    .d1(q_2_7),
    .q(q_3_7)
  );
  

  flop_with_mux u_3_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_7),
    .d1(q_2_8),
    .q(q_3_8)
  );
  

  flop_with_mux u_3_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_8),
    .d1(q_2_9),
    .q(q_3_9)
  );
  

  flop_with_mux u_3_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_9),
    .d1(q_2_10),
    .q(q_3_10)
  );
  

  flop_with_mux u_3_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_10),
    .d1(q_2_11),
    .q(q_3_11)
  );
  

  flop_with_mux u_3_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_11),
    .d1(q_2_12),
    .q(q_3_12)
  );
  

  flop_with_mux u_3_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_12),
    .d1(q_2_13),
    .q(q_3_13)
  );
  

  flop_with_mux u_3_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_13),
    .d1(q_2_14),
    .q(q_3_14)
  );
  

  flop_with_mux u_3_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_14),
    .d1(q_2_15),
    .q(q_3_15)
  );
  

  flop_with_mux u_3_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_15),
    .d1(q_2_16),
    .q(q_3_16)
  );
  

  flop_with_mux u_3_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_16),
    .d1(q_2_17),
    .q(q_3_17)
  );
  

  flop_with_mux u_3_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_17),
    .d1(q_2_18),
    .q(q_3_18)
  );
  

  flop_with_mux u_3_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_18),
    .d1(q_2_19),
    .q(q_3_19)
  );
  

  flop_with_mux u_3_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_19),
    .d1(q_2_20),
    .q(q_3_20)
  );
  

  flop_with_mux u_3_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_20),
    .d1(q_2_21),
    .q(q_3_21)
  );
  

  flop_with_mux u_3_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_21),
    .d1(q_2_22),
    .q(q_3_22)
  );
  

  flop_with_mux u_3_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_22),
    .d1(q_2_23),
    .q(q_3_23)
  );
  

  flop_with_mux u_3_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_23),
    .d1(q_2_24),
    .q(q_3_24)
  );
  

  flop_with_mux u_3_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_24),
    .d1(q_2_25),
    .q(q_3_25)
  );
  

  flop_with_mux u_3_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_25),
    .d1(q_2_26),
    .q(q_3_26)
  );
  

  flop_with_mux u_3_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_26),
    .d1(q_2_27),
    .q(q_3_27)
  );
  

  flop_with_mux u_3_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_27),
    .d1(q_2_28),
    .q(q_3_28)
  );
  

  flop_with_mux u_3_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_28),
    .d1(q_2_29),
    .q(q_3_29)
  );
  

  flop_with_mux u_3_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_29),
    .d1(q_2_30),
    .q(q_3_30)
  );
  

  flop_with_mux u_3_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_30),
    .d1(q_2_31),
    .q(q_3_31)
  );
  

  flop_with_mux u_3_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_31),
    .d1(q_2_32),
    .q(q_3_32)
  );
  

  flop_with_mux u_3_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_32),
    .d1(q_2_33),
    .q(q_3_33)
  );
  

  flop_with_mux u_3_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_33),
    .d1(q_2_34),
    .q(q_3_34)
  );
  

  flop_with_mux u_3_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_34),
    .d1(q_2_35),
    .q(q_3_35)
  );
  

  flop_with_mux u_3_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_35),
    .d1(q_2_36),
    .q(q_3_36)
  );
  

  flop_with_mux u_3_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_36),
    .d1(q_2_37),
    .q(q_3_37)
  );
  

  flop_with_mux u_3_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_37),
    .d1(q_2_38),
    .q(q_3_38)
  );
  

  flop_with_mux u_3_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_38),
    .d1(q_2_39),
    .q(q_3_39)
  );
  

  flop_with_mux u_4_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_minus1),
    .d1(q_3_0),
    .q(q_4_0)
  );
  

  flop_with_mux u_4_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_0),
    .d1(q_3_1),
    .q(q_4_1)
  );
  

  flop_with_mux u_4_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_1),
    .d1(q_3_2),
    .q(q_4_2)
  );
  

  flop_with_mux u_4_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_2),
    .d1(q_3_3),
    .q(q_4_3)
  );
  

  flop_with_mux u_4_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_3),
    .d1(q_3_4),
    .q(q_4_4)
  );
  

  flop_with_mux u_4_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_4),
    .d1(q_3_5),
    .q(q_4_5)
  );
  

  flop_with_mux u_4_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_5),
    .d1(q_3_6),
    .q(q_4_6)
  );
  

  flop_with_mux u_4_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_6),
    .d1(q_3_7),
    .q(q_4_7)
  );
  

  flop_with_mux u_4_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_7),
    .d1(q_3_8),
    .q(q_4_8)
  );
  

  flop_with_mux u_4_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_8),
    .d1(q_3_9),
    .q(q_4_9)
  );
  

  flop_with_mux u_4_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_9),
    .d1(q_3_10),
    .q(q_4_10)
  );
  

  flop_with_mux u_4_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_10),
    .d1(q_3_11),
    .q(q_4_11)
  );
  

  flop_with_mux u_4_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_11),
    .d1(q_3_12),
    .q(q_4_12)
  );
  

  flop_with_mux u_4_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_12),
    .d1(q_3_13),
    .q(q_4_13)
  );
  

  flop_with_mux u_4_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_13),
    .d1(q_3_14),
    .q(q_4_14)
  );
  

  flop_with_mux u_4_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_14),
    .d1(q_3_15),
    .q(q_4_15)
  );
  

  flop_with_mux u_4_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_15),
    .d1(q_3_16),
    .q(q_4_16)
  );
  

  flop_with_mux u_4_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_16),
    .d1(q_3_17),
    .q(q_4_17)
  );
  

  flop_with_mux u_4_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_17),
    .d1(q_3_18),
    .q(q_4_18)
  );
  

  flop_with_mux u_4_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_18),
    .d1(q_3_19),
    .q(q_4_19)
  );
  

  flop_with_mux u_4_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_19),
    .d1(q_3_20),
    .q(q_4_20)
  );
  

  flop_with_mux u_4_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_20),
    .d1(q_3_21),
    .q(q_4_21)
  );
  

  flop_with_mux u_4_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_21),
    .d1(q_3_22),
    .q(q_4_22)
  );
  

  flop_with_mux u_4_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_22),
    .d1(q_3_23),
    .q(q_4_23)
  );
  

  flop_with_mux u_4_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_23),
    .d1(q_3_24),
    .q(q_4_24)
  );
  

  flop_with_mux u_4_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_24),
    .d1(q_3_25),
    .q(q_4_25)
  );
  

  flop_with_mux u_4_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_25),
    .d1(q_3_26),
    .q(q_4_26)
  );
  

  flop_with_mux u_4_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_26),
    .d1(q_3_27),
    .q(q_4_27)
  );
  

  flop_with_mux u_4_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_27),
    .d1(q_3_28),
    .q(q_4_28)
  );
  

  flop_with_mux u_4_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_28),
    .d1(q_3_29),
    .q(q_4_29)
  );
  

  flop_with_mux u_4_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_29),
    .d1(q_3_30),
    .q(q_4_30)
  );
  

  flop_with_mux u_4_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_30),
    .d1(q_3_31),
    .q(q_4_31)
  );
  

  flop_with_mux u_4_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_31),
    .d1(q_3_32),
    .q(q_4_32)
  );
  

  flop_with_mux u_4_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_32),
    .d1(q_3_33),
    .q(q_4_33)
  );
  

  flop_with_mux u_4_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_33),
    .d1(q_3_34),
    .q(q_4_34)
  );
  

  flop_with_mux u_4_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_34),
    .d1(q_3_35),
    .q(q_4_35)
  );
  

  flop_with_mux u_4_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_35),
    .d1(q_3_36),
    .q(q_4_36)
  );
  

  flop_with_mux u_4_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_36),
    .d1(q_3_37),
    .q(q_4_37)
  );
  

  flop_with_mux u_4_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_37),
    .d1(q_3_38),
    .q(q_4_38)
  );
  

  flop_with_mux u_4_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_38),
    .d1(q_3_39),
    .q(q_4_39)
  );
  

  flop_with_mux u_5_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_minus1),
    .d1(q_4_0),
    .q(q_5_0)
  );
  

  flop_with_mux u_5_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_0),
    .d1(q_4_1),
    .q(q_5_1)
  );
  

  flop_with_mux u_5_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_1),
    .d1(q_4_2),
    .q(q_5_2)
  );
  

  flop_with_mux u_5_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_2),
    .d1(q_4_3),
    .q(q_5_3)
  );
  

  flop_with_mux u_5_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_3),
    .d1(q_4_4),
    .q(q_5_4)
  );
  

  flop_with_mux u_5_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_4),
    .d1(q_4_5),
    .q(q_5_5)
  );
  

  flop_with_mux u_5_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_5),
    .d1(q_4_6),
    .q(q_5_6)
  );
  

  flop_with_mux u_5_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_6),
    .d1(q_4_7),
    .q(q_5_7)
  );
  

  flop_with_mux u_5_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_7),
    .d1(q_4_8),
    .q(q_5_8)
  );
  

  flop_with_mux u_5_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_8),
    .d1(q_4_9),
    .q(q_5_9)
  );
  

  flop_with_mux u_5_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_9),
    .d1(q_4_10),
    .q(q_5_10)
  );
  

  flop_with_mux u_5_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_10),
    .d1(q_4_11),
    .q(q_5_11)
  );
  

  flop_with_mux u_5_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_11),
    .d1(q_4_12),
    .q(q_5_12)
  );
  

  flop_with_mux u_5_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_12),
    .d1(q_4_13),
    .q(q_5_13)
  );
  

  flop_with_mux u_5_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_13),
    .d1(q_4_14),
    .q(q_5_14)
  );
  

  flop_with_mux u_5_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_14),
    .d1(q_4_15),
    .q(q_5_15)
  );
  

  flop_with_mux u_5_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_15),
    .d1(q_4_16),
    .q(q_5_16)
  );
  

  flop_with_mux u_5_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_16),
    .d1(q_4_17),
    .q(q_5_17)
  );
  

  flop_with_mux u_5_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_17),
    .d1(q_4_18),
    .q(q_5_18)
  );
  

  flop_with_mux u_5_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_18),
    .d1(q_4_19),
    .q(q_5_19)
  );
  

  flop_with_mux u_5_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_19),
    .d1(q_4_20),
    .q(q_5_20)
  );
  

  flop_with_mux u_5_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_20),
    .d1(q_4_21),
    .q(q_5_21)
  );
  

  flop_with_mux u_5_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_21),
    .d1(q_4_22),
    .q(q_5_22)
  );
  

  flop_with_mux u_5_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_22),
    .d1(q_4_23),
    .q(q_5_23)
  );
  

  flop_with_mux u_5_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_23),
    .d1(q_4_24),
    .q(q_5_24)
  );
  

  flop_with_mux u_5_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_24),
    .d1(q_4_25),
    .q(q_5_25)
  );
  

  flop_with_mux u_5_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_25),
    .d1(q_4_26),
    .q(q_5_26)
  );
  

  flop_with_mux u_5_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_26),
    .d1(q_4_27),
    .q(q_5_27)
  );
  

  flop_with_mux u_5_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_27),
    .d1(q_4_28),
    .q(q_5_28)
  );
  

  flop_with_mux u_5_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_28),
    .d1(q_4_29),
    .q(q_5_29)
  );
  

  flop_with_mux u_5_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_29),
    .d1(q_4_30),
    .q(q_5_30)
  );
  

  flop_with_mux u_5_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_30),
    .d1(q_4_31),
    .q(q_5_31)
  );
  

  flop_with_mux u_5_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_31),
    .d1(q_4_32),
    .q(q_5_32)
  );
  

  flop_with_mux u_5_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_32),
    .d1(q_4_33),
    .q(q_5_33)
  );
  

  flop_with_mux u_5_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_33),
    .d1(q_4_34),
    .q(q_5_34)
  );
  

  flop_with_mux u_5_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_34),
    .d1(q_4_35),
    .q(q_5_35)
  );
  

  flop_with_mux u_5_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_35),
    .d1(q_4_36),
    .q(q_5_36)
  );
  

  flop_with_mux u_5_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_36),
    .d1(q_4_37),
    .q(q_5_37)
  );
  

  flop_with_mux u_5_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_37),
    .d1(q_4_38),
    .q(q_5_38)
  );
  

  flop_with_mux u_5_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_38),
    .d1(q_4_39),
    .q(q_5_39)
  );
  

  flop_with_mux u_6_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_minus1),
    .d1(q_5_0),
    .q(q_6_0)
  );
  

  flop_with_mux u_6_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_0),
    .d1(q_5_1),
    .q(q_6_1)
  );
  

  flop_with_mux u_6_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_1),
    .d1(q_5_2),
    .q(q_6_2)
  );
  

  flop_with_mux u_6_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_2),
    .d1(q_5_3),
    .q(q_6_3)
  );
  

  flop_with_mux u_6_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_3),
    .d1(q_5_4),
    .q(q_6_4)
  );
  

  flop_with_mux u_6_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_4),
    .d1(q_5_5),
    .q(q_6_5)
  );
  

  flop_with_mux u_6_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_5),
    .d1(q_5_6),
    .q(q_6_6)
  );
  

  flop_with_mux u_6_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_6),
    .d1(q_5_7),
    .q(q_6_7)
  );
  

  flop_with_mux u_6_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_7),
    .d1(q_5_8),
    .q(q_6_8)
  );
  

  flop_with_mux u_6_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_8),
    .d1(q_5_9),
    .q(q_6_9)
  );
  

  flop_with_mux u_6_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_9),
    .d1(q_5_10),
    .q(q_6_10)
  );
  

  flop_with_mux u_6_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_10),
    .d1(q_5_11),
    .q(q_6_11)
  );
  

  flop_with_mux u_6_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_11),
    .d1(q_5_12),
    .q(q_6_12)
  );
  

  flop_with_mux u_6_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_12),
    .d1(q_5_13),
    .q(q_6_13)
  );
  

  flop_with_mux u_6_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_13),
    .d1(q_5_14),
    .q(q_6_14)
  );
  

  flop_with_mux u_6_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_14),
    .d1(q_5_15),
    .q(q_6_15)
  );
  

  flop_with_mux u_6_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_15),
    .d1(q_5_16),
    .q(q_6_16)
  );
  

  flop_with_mux u_6_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_16),
    .d1(q_5_17),
    .q(q_6_17)
  );
  

  flop_with_mux u_6_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_17),
    .d1(q_5_18),
    .q(q_6_18)
  );
  

  flop_with_mux u_6_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_18),
    .d1(q_5_19),
    .q(q_6_19)
  );
  

  flop_with_mux u_6_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_19),
    .d1(q_5_20),
    .q(q_6_20)
  );
  

  flop_with_mux u_6_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_20),
    .d1(q_5_21),
    .q(q_6_21)
  );
  

  flop_with_mux u_6_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_21),
    .d1(q_5_22),
    .q(q_6_22)
  );
  

  flop_with_mux u_6_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_22),
    .d1(q_5_23),
    .q(q_6_23)
  );
  

  flop_with_mux u_6_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_23),
    .d1(q_5_24),
    .q(q_6_24)
  );
  

  flop_with_mux u_6_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_24),
    .d1(q_5_25),
    .q(q_6_25)
  );
  

  flop_with_mux u_6_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_25),
    .d1(q_5_26),
    .q(q_6_26)
  );
  

  flop_with_mux u_6_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_26),
    .d1(q_5_27),
    .q(q_6_27)
  );
  

  flop_with_mux u_6_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_27),
    .d1(q_5_28),
    .q(q_6_28)
  );
  

  flop_with_mux u_6_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_28),
    .d1(q_5_29),
    .q(q_6_29)
  );
  

  flop_with_mux u_6_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_29),
    .d1(q_5_30),
    .q(q_6_30)
  );
  

  flop_with_mux u_6_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_30),
    .d1(q_5_31),
    .q(q_6_31)
  );
  

  flop_with_mux u_6_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_31),
    .d1(q_5_32),
    .q(q_6_32)
  );
  

  flop_with_mux u_6_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_32),
    .d1(q_5_33),
    .q(q_6_33)
  );
  

  flop_with_mux u_6_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_33),
    .d1(q_5_34),
    .q(q_6_34)
  );
  

  flop_with_mux u_6_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_34),
    .d1(q_5_35),
    .q(q_6_35)
  );
  

  flop_with_mux u_6_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_35),
    .d1(q_5_36),
    .q(q_6_36)
  );
  

  flop_with_mux u_6_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_36),
    .d1(q_5_37),
    .q(q_6_37)
  );
  

  flop_with_mux u_6_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_37),
    .d1(q_5_38),
    .q(q_6_38)
  );
  

  flop_with_mux u_6_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_38),
    .d1(q_5_39),
    .q(q_6_39)
  );
  

  flop_with_mux u_7_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_minus1),
    .d1(q_6_0),
    .q(q_7_0)
  );
  

  flop_with_mux u_7_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_0),
    .d1(q_6_1),
    .q(q_7_1)
  );
  

  flop_with_mux u_7_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_1),
    .d1(q_6_2),
    .q(q_7_2)
  );
  

  flop_with_mux u_7_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_2),
    .d1(q_6_3),
    .q(q_7_3)
  );
  

  flop_with_mux u_7_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_3),
    .d1(q_6_4),
    .q(q_7_4)
  );
  

  flop_with_mux u_7_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_4),
    .d1(q_6_5),
    .q(q_7_5)
  );
  

  flop_with_mux u_7_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_5),
    .d1(q_6_6),
    .q(q_7_6)
  );
  

  flop_with_mux u_7_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_6),
    .d1(q_6_7),
    .q(q_7_7)
  );
  

  flop_with_mux u_7_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_7),
    .d1(q_6_8),
    .q(q_7_8)
  );
  

  flop_with_mux u_7_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_8),
    .d1(q_6_9),
    .q(q_7_9)
  );
  

  flop_with_mux u_7_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_9),
    .d1(q_6_10),
    .q(q_7_10)
  );
  

  flop_with_mux u_7_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_10),
    .d1(q_6_11),
    .q(q_7_11)
  );
  

  flop_with_mux u_7_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_11),
    .d1(q_6_12),
    .q(q_7_12)
  );
  

  flop_with_mux u_7_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_12),
    .d1(q_6_13),
    .q(q_7_13)
  );
  

  flop_with_mux u_7_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_13),
    .d1(q_6_14),
    .q(q_7_14)
  );
  

  flop_with_mux u_7_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_14),
    .d1(q_6_15),
    .q(q_7_15)
  );
  

  flop_with_mux u_7_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_15),
    .d1(q_6_16),
    .q(q_7_16)
  );
  

  flop_with_mux u_7_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_16),
    .d1(q_6_17),
    .q(q_7_17)
  );
  

  flop_with_mux u_7_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_17),
    .d1(q_6_18),
    .q(q_7_18)
  );
  

  flop_with_mux u_7_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_18),
    .d1(q_6_19),
    .q(q_7_19)
  );
  

  flop_with_mux u_7_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_19),
    .d1(q_6_20),
    .q(q_7_20)
  );
  

  flop_with_mux u_7_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_20),
    .d1(q_6_21),
    .q(q_7_21)
  );
  

  flop_with_mux u_7_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_21),
    .d1(q_6_22),
    .q(q_7_22)
  );
  

  flop_with_mux u_7_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_22),
    .d1(q_6_23),
    .q(q_7_23)
  );
  

  flop_with_mux u_7_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_23),
    .d1(q_6_24),
    .q(q_7_24)
  );
  

  flop_with_mux u_7_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_24),
    .d1(q_6_25),
    .q(q_7_25)
  );
  

  flop_with_mux u_7_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_25),
    .d1(q_6_26),
    .q(q_7_26)
  );
  

  flop_with_mux u_7_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_26),
    .d1(q_6_27),
    .q(q_7_27)
  );
  

  flop_with_mux u_7_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_27),
    .d1(q_6_28),
    .q(q_7_28)
  );
  

  flop_with_mux u_7_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_28),
    .d1(q_6_29),
    .q(q_7_29)
  );
  

  flop_with_mux u_7_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_29),
    .d1(q_6_30),
    .q(q_7_30)
  );
  

  flop_with_mux u_7_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_30),
    .d1(q_6_31),
    .q(q_7_31)
  );
  

  flop_with_mux u_7_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_31),
    .d1(q_6_32),
    .q(q_7_32)
  );
  

  flop_with_mux u_7_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_32),
    .d1(q_6_33),
    .q(q_7_33)
  );
  

  flop_with_mux u_7_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_33),
    .d1(q_6_34),
    .q(q_7_34)
  );
  

  flop_with_mux u_7_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_34),
    .d1(q_6_35),
    .q(q_7_35)
  );
  

  flop_with_mux u_7_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_35),
    .d1(q_6_36),
    .q(q_7_36)
  );
  

  flop_with_mux u_7_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_36),
    .d1(q_6_37),
    .q(q_7_37)
  );
  

  flop_with_mux u_7_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_37),
    .d1(q_6_38),
    .q(q_7_38)
  );
  

  flop_with_mux u_7_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_38),
    .d1(q_6_39),
    .q(q_7_39)
  );
  

  flop_with_mux u_8_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_minus1),
    .d1(q_7_0),
    .q(q_8_0)
  );
  

  flop_with_mux u_8_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_0),
    .d1(q_7_1),
    .q(q_8_1)
  );
  

  flop_with_mux u_8_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_1),
    .d1(q_7_2),
    .q(q_8_2)
  );
  

  flop_with_mux u_8_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_2),
    .d1(q_7_3),
    .q(q_8_3)
  );
  

  flop_with_mux u_8_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_3),
    .d1(q_7_4),
    .q(q_8_4)
  );
  

  flop_with_mux u_8_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_4),
    .d1(q_7_5),
    .q(q_8_5)
  );
  

  flop_with_mux u_8_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_5),
    .d1(q_7_6),
    .q(q_8_6)
  );
  

  flop_with_mux u_8_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_6),
    .d1(q_7_7),
    .q(q_8_7)
  );
  

  flop_with_mux u_8_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_7),
    .d1(q_7_8),
    .q(q_8_8)
  );
  

  flop_with_mux u_8_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_8),
    .d1(q_7_9),
    .q(q_8_9)
  );
  

  flop_with_mux u_8_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_9),
    .d1(q_7_10),
    .q(q_8_10)
  );
  

  flop_with_mux u_8_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_10),
    .d1(q_7_11),
    .q(q_8_11)
  );
  

  flop_with_mux u_8_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_11),
    .d1(q_7_12),
    .q(q_8_12)
  );
  

  flop_with_mux u_8_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_12),
    .d1(q_7_13),
    .q(q_8_13)
  );
  

  flop_with_mux u_8_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_13),
    .d1(q_7_14),
    .q(q_8_14)
  );
  

  flop_with_mux u_8_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_14),
    .d1(q_7_15),
    .q(q_8_15)
  );
  

  flop_with_mux u_8_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_15),
    .d1(q_7_16),
    .q(q_8_16)
  );
  

  flop_with_mux u_8_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_16),
    .d1(q_7_17),
    .q(q_8_17)
  );
  

  flop_with_mux u_8_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_17),
    .d1(q_7_18),
    .q(q_8_18)
  );
  

  flop_with_mux u_8_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_18),
    .d1(q_7_19),
    .q(q_8_19)
  );
  

  flop_with_mux u_8_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_19),
    .d1(q_7_20),
    .q(q_8_20)
  );
  

  flop_with_mux u_8_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_20),
    .d1(q_7_21),
    .q(q_8_21)
  );
  

  flop_with_mux u_8_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_21),
    .d1(q_7_22),
    .q(q_8_22)
  );
  

  flop_with_mux u_8_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_22),
    .d1(q_7_23),
    .q(q_8_23)
  );
  

  flop_with_mux u_8_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_23),
    .d1(q_7_24),
    .q(q_8_24)
  );
  

  flop_with_mux u_8_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_24),
    .d1(q_7_25),
    .q(q_8_25)
  );
  

  flop_with_mux u_8_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_25),
    .d1(q_7_26),
    .q(q_8_26)
  );
  

  flop_with_mux u_8_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_26),
    .d1(q_7_27),
    .q(q_8_27)
  );
  

  flop_with_mux u_8_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_27),
    .d1(q_7_28),
    .q(q_8_28)
  );
  

  flop_with_mux u_8_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_28),
    .d1(q_7_29),
    .q(q_8_29)
  );
  

  flop_with_mux u_8_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_29),
    .d1(q_7_30),
    .q(q_8_30)
  );
  

  flop_with_mux u_8_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_30),
    .d1(q_7_31),
    .q(q_8_31)
  );
  

  flop_with_mux u_8_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_31),
    .d1(q_7_32),
    .q(q_8_32)
  );
  

  flop_with_mux u_8_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_32),
    .d1(q_7_33),
    .q(q_8_33)
  );
  

  flop_with_mux u_8_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_33),
    .d1(q_7_34),
    .q(q_8_34)
  );
  

  flop_with_mux u_8_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_34),
    .d1(q_7_35),
    .q(q_8_35)
  );
  

  flop_with_mux u_8_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_35),
    .d1(q_7_36),
    .q(q_8_36)
  );
  

  flop_with_mux u_8_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_36),
    .d1(q_7_37),
    .q(q_8_37)
  );
  

  flop_with_mux u_8_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_37),
    .d1(q_7_38),
    .q(q_8_38)
  );
  

  flop_with_mux u_8_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_38),
    .d1(q_7_39),
    .q(q_8_39)
  );
  

  flop_with_mux u_9_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_minus1),
    .d1(q_8_0),
    .q(q_9_0)
  );
  

  flop_with_mux u_9_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_0),
    .d1(q_8_1),
    .q(q_9_1)
  );
  

  flop_with_mux u_9_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_1),
    .d1(q_8_2),
    .q(q_9_2)
  );
  

  flop_with_mux u_9_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_2),
    .d1(q_8_3),
    .q(q_9_3)
  );
  

  flop_with_mux u_9_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_3),
    .d1(q_8_4),
    .q(q_9_4)
  );
  

  flop_with_mux u_9_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_4),
    .d1(q_8_5),
    .q(q_9_5)
  );
  

  flop_with_mux u_9_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_5),
    .d1(q_8_6),
    .q(q_9_6)
  );
  

  flop_with_mux u_9_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_6),
    .d1(q_8_7),
    .q(q_9_7)
  );
  

  flop_with_mux u_9_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_7),
    .d1(q_8_8),
    .q(q_9_8)
  );
  

  flop_with_mux u_9_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_8),
    .d1(q_8_9),
    .q(q_9_9)
  );
  

  flop_with_mux u_9_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_9),
    .d1(q_8_10),
    .q(q_9_10)
  );
  

  flop_with_mux u_9_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_10),
    .d1(q_8_11),
    .q(q_9_11)
  );
  

  flop_with_mux u_9_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_11),
    .d1(q_8_12),
    .q(q_9_12)
  );
  

  flop_with_mux u_9_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_12),
    .d1(q_8_13),
    .q(q_9_13)
  );
  

  flop_with_mux u_9_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_13),
    .d1(q_8_14),
    .q(q_9_14)
  );
  

  flop_with_mux u_9_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_14),
    .d1(q_8_15),
    .q(q_9_15)
  );
  

  flop_with_mux u_9_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_15),
    .d1(q_8_16),
    .q(q_9_16)
  );
  

  flop_with_mux u_9_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_16),
    .d1(q_8_17),
    .q(q_9_17)
  );
  

  flop_with_mux u_9_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_17),
    .d1(q_8_18),
    .q(q_9_18)
  );
  

  flop_with_mux u_9_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_18),
    .d1(q_8_19),
    .q(q_9_19)
  );
  

  flop_with_mux u_9_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_19),
    .d1(q_8_20),
    .q(q_9_20)
  );
  

  flop_with_mux u_9_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_20),
    .d1(q_8_21),
    .q(q_9_21)
  );
  

  flop_with_mux u_9_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_21),
    .d1(q_8_22),
    .q(q_9_22)
  );
  

  flop_with_mux u_9_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_22),
    .d1(q_8_23),
    .q(q_9_23)
  );
  

  flop_with_mux u_9_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_23),
    .d1(q_8_24),
    .q(q_9_24)
  );
  

  flop_with_mux u_9_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_24),
    .d1(q_8_25),
    .q(q_9_25)
  );
  

  flop_with_mux u_9_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_25),
    .d1(q_8_26),
    .q(q_9_26)
  );
  

  flop_with_mux u_9_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_26),
    .d1(q_8_27),
    .q(q_9_27)
  );
  

  flop_with_mux u_9_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_27),
    .d1(q_8_28),
    .q(q_9_28)
  );
  

  flop_with_mux u_9_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_28),
    .d1(q_8_29),
    .q(q_9_29)
  );
  

  flop_with_mux u_9_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_29),
    .d1(q_8_30),
    .q(q_9_30)
  );
  

  flop_with_mux u_9_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_30),
    .d1(q_8_31),
    .q(q_9_31)
  );
  

  flop_with_mux u_9_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_31),
    .d1(q_8_32),
    .q(q_9_32)
  );
  

  flop_with_mux u_9_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_32),
    .d1(q_8_33),
    .q(q_9_33)
  );
  

  flop_with_mux u_9_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_33),
    .d1(q_8_34),
    .q(q_9_34)
  );
  

  flop_with_mux u_9_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_34),
    .d1(q_8_35),
    .q(q_9_35)
  );
  

  flop_with_mux u_9_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_35),
    .d1(q_8_36),
    .q(q_9_36)
  );
  

  flop_with_mux u_9_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_36),
    .d1(q_8_37),
    .q(q_9_37)
  );
  

  flop_with_mux u_9_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_37),
    .d1(q_8_38),
    .q(q_9_38)
  );
  

  flop_with_mux u_9_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_38),
    .d1(q_8_39),
    .q(q_9_39)
  );
  

  flop_with_mux u_10_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_minus1),
    .d1(q_9_0),
    .q(q_10_0)
  );
  

  flop_with_mux u_10_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_0),
    .d1(q_9_1),
    .q(q_10_1)
  );
  

  flop_with_mux u_10_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_1),
    .d1(q_9_2),
    .q(q_10_2)
  );
  

  flop_with_mux u_10_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_2),
    .d1(q_9_3),
    .q(q_10_3)
  );
  

  flop_with_mux u_10_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_3),
    .d1(q_9_4),
    .q(q_10_4)
  );
  

  flop_with_mux u_10_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_4),
    .d1(q_9_5),
    .q(q_10_5)
  );
  

  flop_with_mux u_10_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_5),
    .d1(q_9_6),
    .q(q_10_6)
  );
  

  flop_with_mux u_10_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_6),
    .d1(q_9_7),
    .q(q_10_7)
  );
  

  flop_with_mux u_10_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_7),
    .d1(q_9_8),
    .q(q_10_8)
  );
  

  flop_with_mux u_10_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_8),
    .d1(q_9_9),
    .q(q_10_9)
  );
  

  flop_with_mux u_10_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_9),
    .d1(q_9_10),
    .q(q_10_10)
  );
  

  flop_with_mux u_10_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_10),
    .d1(q_9_11),
    .q(q_10_11)
  );
  

  flop_with_mux u_10_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_11),
    .d1(q_9_12),
    .q(q_10_12)
  );
  

  flop_with_mux u_10_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_12),
    .d1(q_9_13),
    .q(q_10_13)
  );
  

  flop_with_mux u_10_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_13),
    .d1(q_9_14),
    .q(q_10_14)
  );
  

  flop_with_mux u_10_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_14),
    .d1(q_9_15),
    .q(q_10_15)
  );
  

  flop_with_mux u_10_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_15),
    .d1(q_9_16),
    .q(q_10_16)
  );
  

  flop_with_mux u_10_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_16),
    .d1(q_9_17),
    .q(q_10_17)
  );
  

  flop_with_mux u_10_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_17),
    .d1(q_9_18),
    .q(q_10_18)
  );
  

  flop_with_mux u_10_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_18),
    .d1(q_9_19),
    .q(q_10_19)
  );
  

  flop_with_mux u_10_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_19),
    .d1(q_9_20),
    .q(q_10_20)
  );
  

  flop_with_mux u_10_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_20),
    .d1(q_9_21),
    .q(q_10_21)
  );
  

  flop_with_mux u_10_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_21),
    .d1(q_9_22),
    .q(q_10_22)
  );
  

  flop_with_mux u_10_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_22),
    .d1(q_9_23),
    .q(q_10_23)
  );
  

  flop_with_mux u_10_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_23),
    .d1(q_9_24),
    .q(q_10_24)
  );
  

  flop_with_mux u_10_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_24),
    .d1(q_9_25),
    .q(q_10_25)
  );
  

  flop_with_mux u_10_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_25),
    .d1(q_9_26),
    .q(q_10_26)
  );
  

  flop_with_mux u_10_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_26),
    .d1(q_9_27),
    .q(q_10_27)
  );
  

  flop_with_mux u_10_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_27),
    .d1(q_9_28),
    .q(q_10_28)
  );
  

  flop_with_mux u_10_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_28),
    .d1(q_9_29),
    .q(q_10_29)
  );
  

  flop_with_mux u_10_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_29),
    .d1(q_9_30),
    .q(q_10_30)
  );
  

  flop_with_mux u_10_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_30),
    .d1(q_9_31),
    .q(q_10_31)
  );
  

  flop_with_mux u_10_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_31),
    .d1(q_9_32),
    .q(q_10_32)
  );
  

  flop_with_mux u_10_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_32),
    .d1(q_9_33),
    .q(q_10_33)
  );
  

  flop_with_mux u_10_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_33),
    .d1(q_9_34),
    .q(q_10_34)
  );
  

  flop_with_mux u_10_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_34),
    .d1(q_9_35),
    .q(q_10_35)
  );
  

  flop_with_mux u_10_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_35),
    .d1(q_9_36),
    .q(q_10_36)
  );
  

  flop_with_mux u_10_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_36),
    .d1(q_9_37),
    .q(q_10_37)
  );
  

  flop_with_mux u_10_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_37),
    .d1(q_9_38),
    .q(q_10_38)
  );
  

  flop_with_mux u_10_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_38),
    .d1(q_9_39),
    .q(q_10_39)
  );
  

  flop_with_mux u_11_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_minus1),
    .d1(q_10_0),
    .q(q_11_0)
  );
  

  flop_with_mux u_11_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_0),
    .d1(q_10_1),
    .q(q_11_1)
  );
  

  flop_with_mux u_11_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_1),
    .d1(q_10_2),
    .q(q_11_2)
  );
  

  flop_with_mux u_11_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_2),
    .d1(q_10_3),
    .q(q_11_3)
  );
  

  flop_with_mux u_11_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_3),
    .d1(q_10_4),
    .q(q_11_4)
  );
  

  flop_with_mux u_11_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_4),
    .d1(q_10_5),
    .q(q_11_5)
  );
  

  flop_with_mux u_11_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_5),
    .d1(q_10_6),
    .q(q_11_6)
  );
  

  flop_with_mux u_11_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_6),
    .d1(q_10_7),
    .q(q_11_7)
  );
  

  flop_with_mux u_11_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_7),
    .d1(q_10_8),
    .q(q_11_8)
  );
  

  flop_with_mux u_11_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_8),
    .d1(q_10_9),
    .q(q_11_9)
  );
  

  flop_with_mux u_11_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_9),
    .d1(q_10_10),
    .q(q_11_10)
  );
  

  flop_with_mux u_11_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_10),
    .d1(q_10_11),
    .q(q_11_11)
  );
  

  flop_with_mux u_11_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_11),
    .d1(q_10_12),
    .q(q_11_12)
  );
  

  flop_with_mux u_11_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_12),
    .d1(q_10_13),
    .q(q_11_13)
  );
  

  flop_with_mux u_11_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_13),
    .d1(q_10_14),
    .q(q_11_14)
  );
  

  flop_with_mux u_11_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_14),
    .d1(q_10_15),
    .q(q_11_15)
  );
  

  flop_with_mux u_11_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_15),
    .d1(q_10_16),
    .q(q_11_16)
  );
  

  flop_with_mux u_11_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_16),
    .d1(q_10_17),
    .q(q_11_17)
  );
  

  flop_with_mux u_11_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_17),
    .d1(q_10_18),
    .q(q_11_18)
  );
  

  flop_with_mux u_11_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_18),
    .d1(q_10_19),
    .q(q_11_19)
  );
  

  flop_with_mux u_11_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_19),
    .d1(q_10_20),
    .q(q_11_20)
  );
  

  flop_with_mux u_11_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_20),
    .d1(q_10_21),
    .q(q_11_21)
  );
  

  flop_with_mux u_11_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_21),
    .d1(q_10_22),
    .q(q_11_22)
  );
  

  flop_with_mux u_11_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_22),
    .d1(q_10_23),
    .q(q_11_23)
  );
  

  flop_with_mux u_11_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_23),
    .d1(q_10_24),
    .q(q_11_24)
  );
  

  flop_with_mux u_11_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_24),
    .d1(q_10_25),
    .q(q_11_25)
  );
  

  flop_with_mux u_11_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_25),
    .d1(q_10_26),
    .q(q_11_26)
  );
  

  flop_with_mux u_11_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_26),
    .d1(q_10_27),
    .q(q_11_27)
  );
  

  flop_with_mux u_11_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_27),
    .d1(q_10_28),
    .q(q_11_28)
  );
  

  flop_with_mux u_11_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_28),
    .d1(q_10_29),
    .q(q_11_29)
  );
  

  flop_with_mux u_11_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_29),
    .d1(q_10_30),
    .q(q_11_30)
  );
  

  flop_with_mux u_11_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_30),
    .d1(q_10_31),
    .q(q_11_31)
  );
  

  flop_with_mux u_11_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_31),
    .d1(q_10_32),
    .q(q_11_32)
  );
  

  flop_with_mux u_11_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_32),
    .d1(q_10_33),
    .q(q_11_33)
  );
  

  flop_with_mux u_11_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_33),
    .d1(q_10_34),
    .q(q_11_34)
  );
  

  flop_with_mux u_11_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_34),
    .d1(q_10_35),
    .q(q_11_35)
  );
  

  flop_with_mux u_11_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_35),
    .d1(q_10_36),
    .q(q_11_36)
  );
  

  flop_with_mux u_11_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_36),
    .d1(q_10_37),
    .q(q_11_37)
  );
  

  flop_with_mux u_11_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_37),
    .d1(q_10_38),
    .q(q_11_38)
  );
  

  flop_with_mux u_11_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_38),
    .d1(q_10_39),
    .q(q_11_39)
  );
  

  flop_with_mux u_12_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_minus1),
    .d1(q_11_0),
    .q(q_12_0)
  );
  

  flop_with_mux u_12_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_0),
    .d1(q_11_1),
    .q(q_12_1)
  );
  

  flop_with_mux u_12_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_1),
    .d1(q_11_2),
    .q(q_12_2)
  );
  

  flop_with_mux u_12_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_2),
    .d1(q_11_3),
    .q(q_12_3)
  );
  

  flop_with_mux u_12_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_3),
    .d1(q_11_4),
    .q(q_12_4)
  );
  

  flop_with_mux u_12_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_4),
    .d1(q_11_5),
    .q(q_12_5)
  );
  

  flop_with_mux u_12_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_5),
    .d1(q_11_6),
    .q(q_12_6)
  );
  

  flop_with_mux u_12_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_6),
    .d1(q_11_7),
    .q(q_12_7)
  );
  

  flop_with_mux u_12_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_7),
    .d1(q_11_8),
    .q(q_12_8)
  );
  

  flop_with_mux u_12_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_8),
    .d1(q_11_9),
    .q(q_12_9)
  );
  

  flop_with_mux u_12_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_9),
    .d1(q_11_10),
    .q(q_12_10)
  );
  

  flop_with_mux u_12_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_10),
    .d1(q_11_11),
    .q(q_12_11)
  );
  

  flop_with_mux u_12_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_11),
    .d1(q_11_12),
    .q(q_12_12)
  );
  

  flop_with_mux u_12_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_12),
    .d1(q_11_13),
    .q(q_12_13)
  );
  

  flop_with_mux u_12_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_13),
    .d1(q_11_14),
    .q(q_12_14)
  );
  

  flop_with_mux u_12_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_14),
    .d1(q_11_15),
    .q(q_12_15)
  );
  

  flop_with_mux u_12_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_15),
    .d1(q_11_16),
    .q(q_12_16)
  );
  

  flop_with_mux u_12_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_16),
    .d1(q_11_17),
    .q(q_12_17)
  );
  

  flop_with_mux u_12_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_17),
    .d1(q_11_18),
    .q(q_12_18)
  );
  

  flop_with_mux u_12_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_18),
    .d1(q_11_19),
    .q(q_12_19)
  );
  

  flop_with_mux u_12_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_19),
    .d1(q_11_20),
    .q(q_12_20)
  );
  

  flop_with_mux u_12_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_20),
    .d1(q_11_21),
    .q(q_12_21)
  );
  

  flop_with_mux u_12_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_21),
    .d1(q_11_22),
    .q(q_12_22)
  );
  

  flop_with_mux u_12_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_22),
    .d1(q_11_23),
    .q(q_12_23)
  );
  

  flop_with_mux u_12_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_23),
    .d1(q_11_24),
    .q(q_12_24)
  );
  

  flop_with_mux u_12_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_24),
    .d1(q_11_25),
    .q(q_12_25)
  );
  

  flop_with_mux u_12_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_25),
    .d1(q_11_26),
    .q(q_12_26)
  );
  

  flop_with_mux u_12_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_26),
    .d1(q_11_27),
    .q(q_12_27)
  );
  

  flop_with_mux u_12_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_27),
    .d1(q_11_28),
    .q(q_12_28)
  );
  

  flop_with_mux u_12_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_28),
    .d1(q_11_29),
    .q(q_12_29)
  );
  

  flop_with_mux u_12_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_29),
    .d1(q_11_30),
    .q(q_12_30)
  );
  

  flop_with_mux u_12_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_30),
    .d1(q_11_31),
    .q(q_12_31)
  );
  

  flop_with_mux u_12_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_31),
    .d1(q_11_32),
    .q(q_12_32)
  );
  

  flop_with_mux u_12_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_32),
    .d1(q_11_33),
    .q(q_12_33)
  );
  

  flop_with_mux u_12_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_33),
    .d1(q_11_34),
    .q(q_12_34)
  );
  

  flop_with_mux u_12_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_34),
    .d1(q_11_35),
    .q(q_12_35)
  );
  

  flop_with_mux u_12_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_35),
    .d1(q_11_36),
    .q(q_12_36)
  );
  

  flop_with_mux u_12_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_36),
    .d1(q_11_37),
    .q(q_12_37)
  );
  

  flop_with_mux u_12_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_37),
    .d1(q_11_38),
    .q(q_12_38)
  );
  

  flop_with_mux u_12_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_38),
    .d1(q_11_39),
    .q(q_12_39)
  );
  

  flop_with_mux u_13_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_minus1),
    .d1(q_12_0),
    .q(q_13_0)
  );
  

  flop_with_mux u_13_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_0),
    .d1(q_12_1),
    .q(q_13_1)
  );
  

  flop_with_mux u_13_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_1),
    .d1(q_12_2),
    .q(q_13_2)
  );
  

  flop_with_mux u_13_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_2),
    .d1(q_12_3),
    .q(q_13_3)
  );
  

  flop_with_mux u_13_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_3),
    .d1(q_12_4),
    .q(q_13_4)
  );
  

  flop_with_mux u_13_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_4),
    .d1(q_12_5),
    .q(q_13_5)
  );
  

  flop_with_mux u_13_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_5),
    .d1(q_12_6),
    .q(q_13_6)
  );
  

  flop_with_mux u_13_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_6),
    .d1(q_12_7),
    .q(q_13_7)
  );
  

  flop_with_mux u_13_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_7),
    .d1(q_12_8),
    .q(q_13_8)
  );
  

  flop_with_mux u_13_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_8),
    .d1(q_12_9),
    .q(q_13_9)
  );
  

  flop_with_mux u_13_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_9),
    .d1(q_12_10),
    .q(q_13_10)
  );
  

  flop_with_mux u_13_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_10),
    .d1(q_12_11),
    .q(q_13_11)
  );
  

  flop_with_mux u_13_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_11),
    .d1(q_12_12),
    .q(q_13_12)
  );
  

  flop_with_mux u_13_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_12),
    .d1(q_12_13),
    .q(q_13_13)
  );
  

  flop_with_mux u_13_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_13),
    .d1(q_12_14),
    .q(q_13_14)
  );
  

  flop_with_mux u_13_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_14),
    .d1(q_12_15),
    .q(q_13_15)
  );
  

  flop_with_mux u_13_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_15),
    .d1(q_12_16),
    .q(q_13_16)
  );
  

  flop_with_mux u_13_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_16),
    .d1(q_12_17),
    .q(q_13_17)
  );
  

  flop_with_mux u_13_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_17),
    .d1(q_12_18),
    .q(q_13_18)
  );
  

  flop_with_mux u_13_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_18),
    .d1(q_12_19),
    .q(q_13_19)
  );
  

  flop_with_mux u_13_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_19),
    .d1(q_12_20),
    .q(q_13_20)
  );
  

  flop_with_mux u_13_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_20),
    .d1(q_12_21),
    .q(q_13_21)
  );
  

  flop_with_mux u_13_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_21),
    .d1(q_12_22),
    .q(q_13_22)
  );
  

  flop_with_mux u_13_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_22),
    .d1(q_12_23),
    .q(q_13_23)
  );
  

  flop_with_mux u_13_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_23),
    .d1(q_12_24),
    .q(q_13_24)
  );
  

  flop_with_mux u_13_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_24),
    .d1(q_12_25),
    .q(q_13_25)
  );
  

  flop_with_mux u_13_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_25),
    .d1(q_12_26),
    .q(q_13_26)
  );
  

  flop_with_mux u_13_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_26),
    .d1(q_12_27),
    .q(q_13_27)
  );
  

  flop_with_mux u_13_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_27),
    .d1(q_12_28),
    .q(q_13_28)
  );
  

  flop_with_mux u_13_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_28),
    .d1(q_12_29),
    .q(q_13_29)
  );
  

  flop_with_mux u_13_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_29),
    .d1(q_12_30),
    .q(q_13_30)
  );
  

  flop_with_mux u_13_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_30),
    .d1(q_12_31),
    .q(q_13_31)
  );
  

  flop_with_mux u_13_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_31),
    .d1(q_12_32),
    .q(q_13_32)
  );
  

  flop_with_mux u_13_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_32),
    .d1(q_12_33),
    .q(q_13_33)
  );
  

  flop_with_mux u_13_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_33),
    .d1(q_12_34),
    .q(q_13_34)
  );
  

  flop_with_mux u_13_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_34),
    .d1(q_12_35),
    .q(q_13_35)
  );
  

  flop_with_mux u_13_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_35),
    .d1(q_12_36),
    .q(q_13_36)
  );
  

  flop_with_mux u_13_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_36),
    .d1(q_12_37),
    .q(q_13_37)
  );
  

  flop_with_mux u_13_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_37),
    .d1(q_12_38),
    .q(q_13_38)
  );
  

  flop_with_mux u_13_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_38),
    .d1(q_12_39),
    .q(q_13_39)
  );
  

  flop_with_mux u_14_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_minus1),
    .d1(q_13_0),
    .q(q_14_0)
  );
  

  flop_with_mux u_14_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_0),
    .d1(q_13_1),
    .q(q_14_1)
  );
  

  flop_with_mux u_14_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_1),
    .d1(q_13_2),
    .q(q_14_2)
  );
  

  flop_with_mux u_14_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_2),
    .d1(q_13_3),
    .q(q_14_3)
  );
  

  flop_with_mux u_14_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_3),
    .d1(q_13_4),
    .q(q_14_4)
  );
  

  flop_with_mux u_14_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_4),
    .d1(q_13_5),
    .q(q_14_5)
  );
  

  flop_with_mux u_14_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_5),
    .d1(q_13_6),
    .q(q_14_6)
  );
  

  flop_with_mux u_14_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_6),
    .d1(q_13_7),
    .q(q_14_7)
  );
  

  flop_with_mux u_14_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_7),
    .d1(q_13_8),
    .q(q_14_8)
  );
  

  flop_with_mux u_14_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_8),
    .d1(q_13_9),
    .q(q_14_9)
  );
  

  flop_with_mux u_14_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_9),
    .d1(q_13_10),
    .q(q_14_10)
  );
  

  flop_with_mux u_14_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_10),
    .d1(q_13_11),
    .q(q_14_11)
  );
  

  flop_with_mux u_14_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_11),
    .d1(q_13_12),
    .q(q_14_12)
  );
  

  flop_with_mux u_14_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_12),
    .d1(q_13_13),
    .q(q_14_13)
  );
  

  flop_with_mux u_14_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_13),
    .d1(q_13_14),
    .q(q_14_14)
  );
  

  flop_with_mux u_14_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_14),
    .d1(q_13_15),
    .q(q_14_15)
  );
  

  flop_with_mux u_14_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_15),
    .d1(q_13_16),
    .q(q_14_16)
  );
  

  flop_with_mux u_14_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_16),
    .d1(q_13_17),
    .q(q_14_17)
  );
  

  flop_with_mux u_14_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_17),
    .d1(q_13_18),
    .q(q_14_18)
  );
  

  flop_with_mux u_14_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_18),
    .d1(q_13_19),
    .q(q_14_19)
  );
  

  flop_with_mux u_14_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_19),
    .d1(q_13_20),
    .q(q_14_20)
  );
  

  flop_with_mux u_14_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_20),
    .d1(q_13_21),
    .q(q_14_21)
  );
  

  flop_with_mux u_14_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_21),
    .d1(q_13_22),
    .q(q_14_22)
  );
  

  flop_with_mux u_14_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_22),
    .d1(q_13_23),
    .q(q_14_23)
  );
  

  flop_with_mux u_14_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_23),
    .d1(q_13_24),
    .q(q_14_24)
  );
  

  flop_with_mux u_14_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_24),
    .d1(q_13_25),
    .q(q_14_25)
  );
  

  flop_with_mux u_14_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_25),
    .d1(q_13_26),
    .q(q_14_26)
  );
  

  flop_with_mux u_14_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_26),
    .d1(q_13_27),
    .q(q_14_27)
  );
  

  flop_with_mux u_14_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_27),
    .d1(q_13_28),
    .q(q_14_28)
  );
  

  flop_with_mux u_14_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_28),
    .d1(q_13_29),
    .q(q_14_29)
  );
  

  flop_with_mux u_14_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_29),
    .d1(q_13_30),
    .q(q_14_30)
  );
  

  flop_with_mux u_14_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_30),
    .d1(q_13_31),
    .q(q_14_31)
  );
  

  flop_with_mux u_14_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_31),
    .d1(q_13_32),
    .q(q_14_32)
  );
  

  flop_with_mux u_14_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_32),
    .d1(q_13_33),
    .q(q_14_33)
  );
  

  flop_with_mux u_14_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_33),
    .d1(q_13_34),
    .q(q_14_34)
  );
  

  flop_with_mux u_14_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_34),
    .d1(q_13_35),
    .q(q_14_35)
  );
  

  flop_with_mux u_14_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_35),
    .d1(q_13_36),
    .q(q_14_36)
  );
  

  flop_with_mux u_14_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_36),
    .d1(q_13_37),
    .q(q_14_37)
  );
  

  flop_with_mux u_14_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_37),
    .d1(q_13_38),
    .q(q_14_38)
  );
  

  flop_with_mux u_14_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_38),
    .d1(q_13_39),
    .q(q_14_39)
  );
  

  flop_with_mux u_15_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_minus1),
    .d1(q_14_0),
    .q(q_15_0)
  );
  

  flop_with_mux u_15_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_0),
    .d1(q_14_1),
    .q(q_15_1)
  );
  

  flop_with_mux u_15_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_1),
    .d1(q_14_2),
    .q(q_15_2)
  );
  

  flop_with_mux u_15_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_2),
    .d1(q_14_3),
    .q(q_15_3)
  );
  

  flop_with_mux u_15_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_3),
    .d1(q_14_4),
    .q(q_15_4)
  );
  

  flop_with_mux u_15_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_4),
    .d1(q_14_5),
    .q(q_15_5)
  );
  

  flop_with_mux u_15_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_5),
    .d1(q_14_6),
    .q(q_15_6)
  );
  

  flop_with_mux u_15_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_6),
    .d1(q_14_7),
    .q(q_15_7)
  );
  

  flop_with_mux u_15_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_7),
    .d1(q_14_8),
    .q(q_15_8)
  );
  

  flop_with_mux u_15_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_8),
    .d1(q_14_9),
    .q(q_15_9)
  );
  

  flop_with_mux u_15_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_9),
    .d1(q_14_10),
    .q(q_15_10)
  );
  

  flop_with_mux u_15_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_10),
    .d1(q_14_11),
    .q(q_15_11)
  );
  

  flop_with_mux u_15_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_11),
    .d1(q_14_12),
    .q(q_15_12)
  );
  

  flop_with_mux u_15_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_12),
    .d1(q_14_13),
    .q(q_15_13)
  );
  

  flop_with_mux u_15_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_13),
    .d1(q_14_14),
    .q(q_15_14)
  );
  

  flop_with_mux u_15_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_14),
    .d1(q_14_15),
    .q(q_15_15)
  );
  

  flop_with_mux u_15_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_15),
    .d1(q_14_16),
    .q(q_15_16)
  );
  

  flop_with_mux u_15_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_16),
    .d1(q_14_17),
    .q(q_15_17)
  );
  

  flop_with_mux u_15_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_17),
    .d1(q_14_18),
    .q(q_15_18)
  );
  

  flop_with_mux u_15_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_18),
    .d1(q_14_19),
    .q(q_15_19)
  );
  

  flop_with_mux u_15_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_19),
    .d1(q_14_20),
    .q(q_15_20)
  );
  

  flop_with_mux u_15_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_20),
    .d1(q_14_21),
    .q(q_15_21)
  );
  

  flop_with_mux u_15_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_21),
    .d1(q_14_22),
    .q(q_15_22)
  );
  

  flop_with_mux u_15_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_22),
    .d1(q_14_23),
    .q(q_15_23)
  );
  

  flop_with_mux u_15_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_23),
    .d1(q_14_24),
    .q(q_15_24)
  );
  

  flop_with_mux u_15_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_24),
    .d1(q_14_25),
    .q(q_15_25)
  );
  

  flop_with_mux u_15_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_25),
    .d1(q_14_26),
    .q(q_15_26)
  );
  

  flop_with_mux u_15_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_26),
    .d1(q_14_27),
    .q(q_15_27)
  );
  

  flop_with_mux u_15_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_27),
    .d1(q_14_28),
    .q(q_15_28)
  );
  

  flop_with_mux u_15_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_28),
    .d1(q_14_29),
    .q(q_15_29)
  );
  

  flop_with_mux u_15_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_29),
    .d1(q_14_30),
    .q(q_15_30)
  );
  

  flop_with_mux u_15_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_30),
    .d1(q_14_31),
    .q(q_15_31)
  );
  

  flop_with_mux u_15_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_31),
    .d1(q_14_32),
    .q(q_15_32)
  );
  

  flop_with_mux u_15_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_32),
    .d1(q_14_33),
    .q(q_15_33)
  );
  

  flop_with_mux u_15_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_33),
    .d1(q_14_34),
    .q(q_15_34)
  );
  

  flop_with_mux u_15_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_34),
    .d1(q_14_35),
    .q(q_15_35)
  );
  

  flop_with_mux u_15_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_35),
    .d1(q_14_36),
    .q(q_15_36)
  );
  

  flop_with_mux u_15_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_36),
    .d1(q_14_37),
    .q(q_15_37)
  );
  

  flop_with_mux u_15_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_37),
    .d1(q_14_38),
    .q(q_15_38)
  );
  

  flop_with_mux u_15_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_38),
    .d1(q_14_39),
    .q(q_15_39)
  );
  

  flop_with_mux u_16_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_minus1),
    .d1(q_15_0),
    .q(q_16_0)
  );
  

  flop_with_mux u_16_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_0),
    .d1(q_15_1),
    .q(q_16_1)
  );
  

  flop_with_mux u_16_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_1),
    .d1(q_15_2),
    .q(q_16_2)
  );
  

  flop_with_mux u_16_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_2),
    .d1(q_15_3),
    .q(q_16_3)
  );
  

  flop_with_mux u_16_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_3),
    .d1(q_15_4),
    .q(q_16_4)
  );
  

  flop_with_mux u_16_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_4),
    .d1(q_15_5),
    .q(q_16_5)
  );
  

  flop_with_mux u_16_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_5),
    .d1(q_15_6),
    .q(q_16_6)
  );
  

  flop_with_mux u_16_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_6),
    .d1(q_15_7),
    .q(q_16_7)
  );
  

  flop_with_mux u_16_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_7),
    .d1(q_15_8),
    .q(q_16_8)
  );
  

  flop_with_mux u_16_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_8),
    .d1(q_15_9),
    .q(q_16_9)
  );
  

  flop_with_mux u_16_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_9),
    .d1(q_15_10),
    .q(q_16_10)
  );
  

  flop_with_mux u_16_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_10),
    .d1(q_15_11),
    .q(q_16_11)
  );
  

  flop_with_mux u_16_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_11),
    .d1(q_15_12),
    .q(q_16_12)
  );
  

  flop_with_mux u_16_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_12),
    .d1(q_15_13),
    .q(q_16_13)
  );
  

  flop_with_mux u_16_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_13),
    .d1(q_15_14),
    .q(q_16_14)
  );
  

  flop_with_mux u_16_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_14),
    .d1(q_15_15),
    .q(q_16_15)
  );
  

  flop_with_mux u_16_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_15),
    .d1(q_15_16),
    .q(q_16_16)
  );
  

  flop_with_mux u_16_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_16),
    .d1(q_15_17),
    .q(q_16_17)
  );
  

  flop_with_mux u_16_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_17),
    .d1(q_15_18),
    .q(q_16_18)
  );
  

  flop_with_mux u_16_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_18),
    .d1(q_15_19),
    .q(q_16_19)
  );
  

  flop_with_mux u_16_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_19),
    .d1(q_15_20),
    .q(q_16_20)
  );
  

  flop_with_mux u_16_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_20),
    .d1(q_15_21),
    .q(q_16_21)
  );
  

  flop_with_mux u_16_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_21),
    .d1(q_15_22),
    .q(q_16_22)
  );
  

  flop_with_mux u_16_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_22),
    .d1(q_15_23),
    .q(q_16_23)
  );
  

  flop_with_mux u_16_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_23),
    .d1(q_15_24),
    .q(q_16_24)
  );
  

  flop_with_mux u_16_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_24),
    .d1(q_15_25),
    .q(q_16_25)
  );
  

  flop_with_mux u_16_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_25),
    .d1(q_15_26),
    .q(q_16_26)
  );
  

  flop_with_mux u_16_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_26),
    .d1(q_15_27),
    .q(q_16_27)
  );
  

  flop_with_mux u_16_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_27),
    .d1(q_15_28),
    .q(q_16_28)
  );
  

  flop_with_mux u_16_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_28),
    .d1(q_15_29),
    .q(q_16_29)
  );
  

  flop_with_mux u_16_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_29),
    .d1(q_15_30),
    .q(q_16_30)
  );
  

  flop_with_mux u_16_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_30),
    .d1(q_15_31),
    .q(q_16_31)
  );
  

  flop_with_mux u_16_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_31),
    .d1(q_15_32),
    .q(q_16_32)
  );
  

  flop_with_mux u_16_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_32),
    .d1(q_15_33),
    .q(q_16_33)
  );
  

  flop_with_mux u_16_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_33),
    .d1(q_15_34),
    .q(q_16_34)
  );
  

  flop_with_mux u_16_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_34),
    .d1(q_15_35),
    .q(q_16_35)
  );
  

  flop_with_mux u_16_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_35),
    .d1(q_15_36),
    .q(q_16_36)
  );
  

  flop_with_mux u_16_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_36),
    .d1(q_15_37),
    .q(q_16_37)
  );
  

  flop_with_mux u_16_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_37),
    .d1(q_15_38),
    .q(q_16_38)
  );
  

  flop_with_mux u_16_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_38),
    .d1(q_15_39),
    .q(q_16_39)
  );
  

  flop_with_mux u_17_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_minus1),
    .d1(q_16_0),
    .q(q_17_0)
  );
  

  flop_with_mux u_17_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_0),
    .d1(q_16_1),
    .q(q_17_1)
  );
  

  flop_with_mux u_17_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_1),
    .d1(q_16_2),
    .q(q_17_2)
  );
  

  flop_with_mux u_17_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_2),
    .d1(q_16_3),
    .q(q_17_3)
  );
  

  flop_with_mux u_17_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_3),
    .d1(q_16_4),
    .q(q_17_4)
  );
  

  flop_with_mux u_17_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_4),
    .d1(q_16_5),
    .q(q_17_5)
  );
  

  flop_with_mux u_17_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_5),
    .d1(q_16_6),
    .q(q_17_6)
  );
  

  flop_with_mux u_17_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_6),
    .d1(q_16_7),
    .q(q_17_7)
  );
  

  flop_with_mux u_17_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_7),
    .d1(q_16_8),
    .q(q_17_8)
  );
  

  flop_with_mux u_17_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_8),
    .d1(q_16_9),
    .q(q_17_9)
  );
  

  flop_with_mux u_17_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_9),
    .d1(q_16_10),
    .q(q_17_10)
  );
  

  flop_with_mux u_17_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_10),
    .d1(q_16_11),
    .q(q_17_11)
  );
  

  flop_with_mux u_17_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_11),
    .d1(q_16_12),
    .q(q_17_12)
  );
  

  flop_with_mux u_17_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_12),
    .d1(q_16_13),
    .q(q_17_13)
  );
  

  flop_with_mux u_17_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_13),
    .d1(q_16_14),
    .q(q_17_14)
  );
  

  flop_with_mux u_17_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_14),
    .d1(q_16_15),
    .q(q_17_15)
  );
  

  flop_with_mux u_17_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_15),
    .d1(q_16_16),
    .q(q_17_16)
  );
  

  flop_with_mux u_17_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_16),
    .d1(q_16_17),
    .q(q_17_17)
  );
  

  flop_with_mux u_17_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_17),
    .d1(q_16_18),
    .q(q_17_18)
  );
  

  flop_with_mux u_17_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_18),
    .d1(q_16_19),
    .q(q_17_19)
  );
  

  flop_with_mux u_17_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_19),
    .d1(q_16_20),
    .q(q_17_20)
  );
  

  flop_with_mux u_17_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_20),
    .d1(q_16_21),
    .q(q_17_21)
  );
  

  flop_with_mux u_17_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_21),
    .d1(q_16_22),
    .q(q_17_22)
  );
  

  flop_with_mux u_17_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_22),
    .d1(q_16_23),
    .q(q_17_23)
  );
  

  flop_with_mux u_17_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_23),
    .d1(q_16_24),
    .q(q_17_24)
  );
  

  flop_with_mux u_17_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_24),
    .d1(q_16_25),
    .q(q_17_25)
  );
  

  flop_with_mux u_17_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_25),
    .d1(q_16_26),
    .q(q_17_26)
  );
  

  flop_with_mux u_17_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_26),
    .d1(q_16_27),
    .q(q_17_27)
  );
  

  flop_with_mux u_17_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_27),
    .d1(q_16_28),
    .q(q_17_28)
  );
  

  flop_with_mux u_17_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_28),
    .d1(q_16_29),
    .q(q_17_29)
  );
  

  flop_with_mux u_17_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_29),
    .d1(q_16_30),
    .q(q_17_30)
  );
  

  flop_with_mux u_17_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_30),
    .d1(q_16_31),
    .q(q_17_31)
  );
  

  flop_with_mux u_17_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_31),
    .d1(q_16_32),
    .q(q_17_32)
  );
  

  flop_with_mux u_17_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_32),
    .d1(q_16_33),
    .q(q_17_33)
  );
  

  flop_with_mux u_17_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_33),
    .d1(q_16_34),
    .q(q_17_34)
  );
  

  flop_with_mux u_17_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_34),
    .d1(q_16_35),
    .q(q_17_35)
  );
  

  flop_with_mux u_17_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_35),
    .d1(q_16_36),
    .q(q_17_36)
  );
  

  flop_with_mux u_17_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_36),
    .d1(q_16_37),
    .q(q_17_37)
  );
  

  flop_with_mux u_17_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_37),
    .d1(q_16_38),
    .q(q_17_38)
  );
  

  flop_with_mux u_17_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_38),
    .d1(q_16_39),
    .q(q_17_39)
  );
  

  flop_with_mux u_18_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_minus1),
    .d1(q_17_0),
    .q(q_18_0)
  );
  

  flop_with_mux u_18_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_0),
    .d1(q_17_1),
    .q(q_18_1)
  );
  

  flop_with_mux u_18_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_1),
    .d1(q_17_2),
    .q(q_18_2)
  );
  

  flop_with_mux u_18_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_2),
    .d1(q_17_3),
    .q(q_18_3)
  );
  

  flop_with_mux u_18_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_3),
    .d1(q_17_4),
    .q(q_18_4)
  );
  

  flop_with_mux u_18_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_4),
    .d1(q_17_5),
    .q(q_18_5)
  );
  

  flop_with_mux u_18_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_5),
    .d1(q_17_6),
    .q(q_18_6)
  );
  

  flop_with_mux u_18_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_6),
    .d1(q_17_7),
    .q(q_18_7)
  );
  

  flop_with_mux u_18_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_7),
    .d1(q_17_8),
    .q(q_18_8)
  );
  

  flop_with_mux u_18_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_8),
    .d1(q_17_9),
    .q(q_18_9)
  );
  

  flop_with_mux u_18_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_9),
    .d1(q_17_10),
    .q(q_18_10)
  );
  

  flop_with_mux u_18_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_10),
    .d1(q_17_11),
    .q(q_18_11)
  );
  

  flop_with_mux u_18_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_11),
    .d1(q_17_12),
    .q(q_18_12)
  );
  

  flop_with_mux u_18_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_12),
    .d1(q_17_13),
    .q(q_18_13)
  );
  

  flop_with_mux u_18_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_13),
    .d1(q_17_14),
    .q(q_18_14)
  );
  

  flop_with_mux u_18_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_14),
    .d1(q_17_15),
    .q(q_18_15)
  );
  

  flop_with_mux u_18_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_15),
    .d1(q_17_16),
    .q(q_18_16)
  );
  

  flop_with_mux u_18_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_16),
    .d1(q_17_17),
    .q(q_18_17)
  );
  

  flop_with_mux u_18_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_17),
    .d1(q_17_18),
    .q(q_18_18)
  );
  

  flop_with_mux u_18_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_18),
    .d1(q_17_19),
    .q(q_18_19)
  );
  

  flop_with_mux u_18_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_19),
    .d1(q_17_20),
    .q(q_18_20)
  );
  

  flop_with_mux u_18_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_20),
    .d1(q_17_21),
    .q(q_18_21)
  );
  

  flop_with_mux u_18_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_21),
    .d1(q_17_22),
    .q(q_18_22)
  );
  

  flop_with_mux u_18_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_22),
    .d1(q_17_23),
    .q(q_18_23)
  );
  

  flop_with_mux u_18_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_23),
    .d1(q_17_24),
    .q(q_18_24)
  );
  

  flop_with_mux u_18_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_24),
    .d1(q_17_25),
    .q(q_18_25)
  );
  

  flop_with_mux u_18_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_25),
    .d1(q_17_26),
    .q(q_18_26)
  );
  

  flop_with_mux u_18_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_26),
    .d1(q_17_27),
    .q(q_18_27)
  );
  

  flop_with_mux u_18_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_27),
    .d1(q_17_28),
    .q(q_18_28)
  );
  

  flop_with_mux u_18_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_28),
    .d1(q_17_29),
    .q(q_18_29)
  );
  

  flop_with_mux u_18_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_29),
    .d1(q_17_30),
    .q(q_18_30)
  );
  

  flop_with_mux u_18_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_30),
    .d1(q_17_31),
    .q(q_18_31)
  );
  

  flop_with_mux u_18_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_31),
    .d1(q_17_32),
    .q(q_18_32)
  );
  

  flop_with_mux u_18_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_32),
    .d1(q_17_33),
    .q(q_18_33)
  );
  

  flop_with_mux u_18_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_33),
    .d1(q_17_34),
    .q(q_18_34)
  );
  

  flop_with_mux u_18_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_34),
    .d1(q_17_35),
    .q(q_18_35)
  );
  

  flop_with_mux u_18_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_35),
    .d1(q_17_36),
    .q(q_18_36)
  );
  

  flop_with_mux u_18_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_36),
    .d1(q_17_37),
    .q(q_18_37)
  );
  

  flop_with_mux u_18_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_37),
    .d1(q_17_38),
    .q(q_18_38)
  );
  

  flop_with_mux u_18_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_38),
    .d1(q_17_39),
    .q(q_18_39)
  );
  

  flop_with_mux u_19_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_minus1),
    .d1(q_18_0),
    .q(q_19_0)
  );
  

  flop_with_mux u_19_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_0),
    .d1(q_18_1),
    .q(q_19_1)
  );
  

  flop_with_mux u_19_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_1),
    .d1(q_18_2),
    .q(q_19_2)
  );
  

  flop_with_mux u_19_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_2),
    .d1(q_18_3),
    .q(q_19_3)
  );
  

  flop_with_mux u_19_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_3),
    .d1(q_18_4),
    .q(q_19_4)
  );
  

  flop_with_mux u_19_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_4),
    .d1(q_18_5),
    .q(q_19_5)
  );
  

  flop_with_mux u_19_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_5),
    .d1(q_18_6),
    .q(q_19_6)
  );
  

  flop_with_mux u_19_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_6),
    .d1(q_18_7),
    .q(q_19_7)
  );
  

  flop_with_mux u_19_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_7),
    .d1(q_18_8),
    .q(q_19_8)
  );
  

  flop_with_mux u_19_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_8),
    .d1(q_18_9),
    .q(q_19_9)
  );
  

  flop_with_mux u_19_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_9),
    .d1(q_18_10),
    .q(q_19_10)
  );
  

  flop_with_mux u_19_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_10),
    .d1(q_18_11),
    .q(q_19_11)
  );
  

  flop_with_mux u_19_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_11),
    .d1(q_18_12),
    .q(q_19_12)
  );
  

  flop_with_mux u_19_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_12),
    .d1(q_18_13),
    .q(q_19_13)
  );
  

  flop_with_mux u_19_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_13),
    .d1(q_18_14),
    .q(q_19_14)
  );
  

  flop_with_mux u_19_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_14),
    .d1(q_18_15),
    .q(q_19_15)
  );
  

  flop_with_mux u_19_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_15),
    .d1(q_18_16),
    .q(q_19_16)
  );
  

  flop_with_mux u_19_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_16),
    .d1(q_18_17),
    .q(q_19_17)
  );
  

  flop_with_mux u_19_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_17),
    .d1(q_18_18),
    .q(q_19_18)
  );
  

  flop_with_mux u_19_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_18),
    .d1(q_18_19),
    .q(q_19_19)
  );
  

  flop_with_mux u_19_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_19),
    .d1(q_18_20),
    .q(q_19_20)
  );
  

  flop_with_mux u_19_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_20),
    .d1(q_18_21),
    .q(q_19_21)
  );
  

  flop_with_mux u_19_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_21),
    .d1(q_18_22),
    .q(q_19_22)
  );
  

  flop_with_mux u_19_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_22),
    .d1(q_18_23),
    .q(q_19_23)
  );
  

  flop_with_mux u_19_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_23),
    .d1(q_18_24),
    .q(q_19_24)
  );
  

  flop_with_mux u_19_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_24),
    .d1(q_18_25),
    .q(q_19_25)
  );
  

  flop_with_mux u_19_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_25),
    .d1(q_18_26),
    .q(q_19_26)
  );
  

  flop_with_mux u_19_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_26),
    .d1(q_18_27),
    .q(q_19_27)
  );
  

  flop_with_mux u_19_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_27),
    .d1(q_18_28),
    .q(q_19_28)
  );
  

  flop_with_mux u_19_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_28),
    .d1(q_18_29),
    .q(q_19_29)
  );
  

  flop_with_mux u_19_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_29),
    .d1(q_18_30),
    .q(q_19_30)
  );
  

  flop_with_mux u_19_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_30),
    .d1(q_18_31),
    .q(q_19_31)
  );
  

  flop_with_mux u_19_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_31),
    .d1(q_18_32),
    .q(q_19_32)
  );
  

  flop_with_mux u_19_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_32),
    .d1(q_18_33),
    .q(q_19_33)
  );
  

  flop_with_mux u_19_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_33),
    .d1(q_18_34),
    .q(q_19_34)
  );
  

  flop_with_mux u_19_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_34),
    .d1(q_18_35),
    .q(q_19_35)
  );
  

  flop_with_mux u_19_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_35),
    .d1(q_18_36),
    .q(q_19_36)
  );
  

  flop_with_mux u_19_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_36),
    .d1(q_18_37),
    .q(q_19_37)
  );
  

  flop_with_mux u_19_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_37),
    .d1(q_18_38),
    .q(q_19_38)
  );
  

  flop_with_mux u_19_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_38),
    .d1(q_18_39),
    .q(q_19_39)
  );
  

  flop_with_mux u_20_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_minus1),
    .d1(q_19_0),
    .q(q_20_0)
  );
  

  flop_with_mux u_20_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_0),
    .d1(q_19_1),
    .q(q_20_1)
  );
  

  flop_with_mux u_20_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_1),
    .d1(q_19_2),
    .q(q_20_2)
  );
  

  flop_with_mux u_20_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_2),
    .d1(q_19_3),
    .q(q_20_3)
  );
  

  flop_with_mux u_20_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_3),
    .d1(q_19_4),
    .q(q_20_4)
  );
  

  flop_with_mux u_20_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_4),
    .d1(q_19_5),
    .q(q_20_5)
  );
  

  flop_with_mux u_20_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_5),
    .d1(q_19_6),
    .q(q_20_6)
  );
  

  flop_with_mux u_20_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_6),
    .d1(q_19_7),
    .q(q_20_7)
  );
  

  flop_with_mux u_20_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_7),
    .d1(q_19_8),
    .q(q_20_8)
  );
  

  flop_with_mux u_20_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_8),
    .d1(q_19_9),
    .q(q_20_9)
  );
  

  flop_with_mux u_20_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_9),
    .d1(q_19_10),
    .q(q_20_10)
  );
  

  flop_with_mux u_20_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_10),
    .d1(q_19_11),
    .q(q_20_11)
  );
  

  flop_with_mux u_20_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_11),
    .d1(q_19_12),
    .q(q_20_12)
  );
  

  flop_with_mux u_20_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_12),
    .d1(q_19_13),
    .q(q_20_13)
  );
  

  flop_with_mux u_20_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_13),
    .d1(q_19_14),
    .q(q_20_14)
  );
  

  flop_with_mux u_20_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_14),
    .d1(q_19_15),
    .q(q_20_15)
  );
  

  flop_with_mux u_20_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_15),
    .d1(q_19_16),
    .q(q_20_16)
  );
  

  flop_with_mux u_20_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_16),
    .d1(q_19_17),
    .q(q_20_17)
  );
  

  flop_with_mux u_20_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_17),
    .d1(q_19_18),
    .q(q_20_18)
  );
  

  flop_with_mux u_20_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_18),
    .d1(q_19_19),
    .q(q_20_19)
  );
  

  flop_with_mux u_20_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_19),
    .d1(q_19_20),
    .q(q_20_20)
  );
  

  flop_with_mux u_20_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_20),
    .d1(q_19_21),
    .q(q_20_21)
  );
  

  flop_with_mux u_20_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_21),
    .d1(q_19_22),
    .q(q_20_22)
  );
  

  flop_with_mux u_20_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_22),
    .d1(q_19_23),
    .q(q_20_23)
  );
  

  flop_with_mux u_20_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_23),
    .d1(q_19_24),
    .q(q_20_24)
  );
  

  flop_with_mux u_20_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_24),
    .d1(q_19_25),
    .q(q_20_25)
  );
  

  flop_with_mux u_20_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_25),
    .d1(q_19_26),
    .q(q_20_26)
  );
  

  flop_with_mux u_20_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_26),
    .d1(q_19_27),
    .q(q_20_27)
  );
  

  flop_with_mux u_20_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_27),
    .d1(q_19_28),
    .q(q_20_28)
  );
  

  flop_with_mux u_20_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_28),
    .d1(q_19_29),
    .q(q_20_29)
  );
  

  flop_with_mux u_20_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_29),
    .d1(q_19_30),
    .q(q_20_30)
  );
  

  flop_with_mux u_20_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_30),
    .d1(q_19_31),
    .q(q_20_31)
  );
  

  flop_with_mux u_20_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_31),
    .d1(q_19_32),
    .q(q_20_32)
  );
  

  flop_with_mux u_20_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_32),
    .d1(q_19_33),
    .q(q_20_33)
  );
  

  flop_with_mux u_20_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_33),
    .d1(q_19_34),
    .q(q_20_34)
  );
  

  flop_with_mux u_20_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_34),
    .d1(q_19_35),
    .q(q_20_35)
  );
  

  flop_with_mux u_20_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_35),
    .d1(q_19_36),
    .q(q_20_36)
  );
  

  flop_with_mux u_20_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_36),
    .d1(q_19_37),
    .q(q_20_37)
  );
  

  flop_with_mux u_20_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_37),
    .d1(q_19_38),
    .q(q_20_38)
  );
  

  flop_with_mux u_20_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_38),
    .d1(q_19_39),
    .q(q_20_39)
  );
  

  flop_with_mux u_21_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_minus1),
    .d1(q_20_0),
    .q(q_21_0)
  );
  

  flop_with_mux u_21_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_0),
    .d1(q_20_1),
    .q(q_21_1)
  );
  

  flop_with_mux u_21_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_1),
    .d1(q_20_2),
    .q(q_21_2)
  );
  

  flop_with_mux u_21_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_2),
    .d1(q_20_3),
    .q(q_21_3)
  );
  

  flop_with_mux u_21_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_3),
    .d1(q_20_4),
    .q(q_21_4)
  );
  

  flop_with_mux u_21_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_4),
    .d1(q_20_5),
    .q(q_21_5)
  );
  

  flop_with_mux u_21_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_5),
    .d1(q_20_6),
    .q(q_21_6)
  );
  

  flop_with_mux u_21_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_6),
    .d1(q_20_7),
    .q(q_21_7)
  );
  

  flop_with_mux u_21_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_7),
    .d1(q_20_8),
    .q(q_21_8)
  );
  

  flop_with_mux u_21_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_8),
    .d1(q_20_9),
    .q(q_21_9)
  );
  

  flop_with_mux u_21_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_9),
    .d1(q_20_10),
    .q(q_21_10)
  );
  

  flop_with_mux u_21_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_10),
    .d1(q_20_11),
    .q(q_21_11)
  );
  

  flop_with_mux u_21_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_11),
    .d1(q_20_12),
    .q(q_21_12)
  );
  

  flop_with_mux u_21_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_12),
    .d1(q_20_13),
    .q(q_21_13)
  );
  

  flop_with_mux u_21_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_13),
    .d1(q_20_14),
    .q(q_21_14)
  );
  

  flop_with_mux u_21_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_14),
    .d1(q_20_15),
    .q(q_21_15)
  );
  

  flop_with_mux u_21_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_15),
    .d1(q_20_16),
    .q(q_21_16)
  );
  

  flop_with_mux u_21_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_16),
    .d1(q_20_17),
    .q(q_21_17)
  );
  

  flop_with_mux u_21_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_17),
    .d1(q_20_18),
    .q(q_21_18)
  );
  

  flop_with_mux u_21_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_18),
    .d1(q_20_19),
    .q(q_21_19)
  );
  

  flop_with_mux u_21_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_19),
    .d1(q_20_20),
    .q(q_21_20)
  );
  

  flop_with_mux u_21_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_20),
    .d1(q_20_21),
    .q(q_21_21)
  );
  

  flop_with_mux u_21_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_21),
    .d1(q_20_22),
    .q(q_21_22)
  );
  

  flop_with_mux u_21_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_22),
    .d1(q_20_23),
    .q(q_21_23)
  );
  

  flop_with_mux u_21_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_23),
    .d1(q_20_24),
    .q(q_21_24)
  );
  

  flop_with_mux u_21_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_24),
    .d1(q_20_25),
    .q(q_21_25)
  );
  

  flop_with_mux u_21_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_25),
    .d1(q_20_26),
    .q(q_21_26)
  );
  

  flop_with_mux u_21_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_26),
    .d1(q_20_27),
    .q(q_21_27)
  );
  

  flop_with_mux u_21_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_27),
    .d1(q_20_28),
    .q(q_21_28)
  );
  

  flop_with_mux u_21_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_28),
    .d1(q_20_29),
    .q(q_21_29)
  );
  

  flop_with_mux u_21_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_29),
    .d1(q_20_30),
    .q(q_21_30)
  );
  

  flop_with_mux u_21_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_30),
    .d1(q_20_31),
    .q(q_21_31)
  );
  

  flop_with_mux u_21_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_31),
    .d1(q_20_32),
    .q(q_21_32)
  );
  

  flop_with_mux u_21_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_32),
    .d1(q_20_33),
    .q(q_21_33)
  );
  

  flop_with_mux u_21_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_33),
    .d1(q_20_34),
    .q(q_21_34)
  );
  

  flop_with_mux u_21_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_34),
    .d1(q_20_35),
    .q(q_21_35)
  );
  

  flop_with_mux u_21_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_35),
    .d1(q_20_36),
    .q(q_21_36)
  );
  

  flop_with_mux u_21_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_36),
    .d1(q_20_37),
    .q(q_21_37)
  );
  

  flop_with_mux u_21_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_37),
    .d1(q_20_38),
    .q(q_21_38)
  );
  

  flop_with_mux u_21_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_38),
    .d1(q_20_39),
    .q(q_21_39)
  );
  

  flop_with_mux u_22_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_minus1),
    .d1(q_21_0),
    .q(q_22_0)
  );
  

  flop_with_mux u_22_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_0),
    .d1(q_21_1),
    .q(q_22_1)
  );
  

  flop_with_mux u_22_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_1),
    .d1(q_21_2),
    .q(q_22_2)
  );
  

  flop_with_mux u_22_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_2),
    .d1(q_21_3),
    .q(q_22_3)
  );
  

  flop_with_mux u_22_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_3),
    .d1(q_21_4),
    .q(q_22_4)
  );
  

  flop_with_mux u_22_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_4),
    .d1(q_21_5),
    .q(q_22_5)
  );
  

  flop_with_mux u_22_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_5),
    .d1(q_21_6),
    .q(q_22_6)
  );
  

  flop_with_mux u_22_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_6),
    .d1(q_21_7),
    .q(q_22_7)
  );
  

  flop_with_mux u_22_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_7),
    .d1(q_21_8),
    .q(q_22_8)
  );
  

  flop_with_mux u_22_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_8),
    .d1(q_21_9),
    .q(q_22_9)
  );
  

  flop_with_mux u_22_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_9),
    .d1(q_21_10),
    .q(q_22_10)
  );
  

  flop_with_mux u_22_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_10),
    .d1(q_21_11),
    .q(q_22_11)
  );
  

  flop_with_mux u_22_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_11),
    .d1(q_21_12),
    .q(q_22_12)
  );
  

  flop_with_mux u_22_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_12),
    .d1(q_21_13),
    .q(q_22_13)
  );
  

  flop_with_mux u_22_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_13),
    .d1(q_21_14),
    .q(q_22_14)
  );
  

  flop_with_mux u_22_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_14),
    .d1(q_21_15),
    .q(q_22_15)
  );
  

  flop_with_mux u_22_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_15),
    .d1(q_21_16),
    .q(q_22_16)
  );
  

  flop_with_mux u_22_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_16),
    .d1(q_21_17),
    .q(q_22_17)
  );
  

  flop_with_mux u_22_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_17),
    .d1(q_21_18),
    .q(q_22_18)
  );
  

  flop_with_mux u_22_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_18),
    .d1(q_21_19),
    .q(q_22_19)
  );
  

  flop_with_mux u_22_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_19),
    .d1(q_21_20),
    .q(q_22_20)
  );
  

  flop_with_mux u_22_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_20),
    .d1(q_21_21),
    .q(q_22_21)
  );
  

  flop_with_mux u_22_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_21),
    .d1(q_21_22),
    .q(q_22_22)
  );
  

  flop_with_mux u_22_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_22),
    .d1(q_21_23),
    .q(q_22_23)
  );
  

  flop_with_mux u_22_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_23),
    .d1(q_21_24),
    .q(q_22_24)
  );
  

  flop_with_mux u_22_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_24),
    .d1(q_21_25),
    .q(q_22_25)
  );
  

  flop_with_mux u_22_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_25),
    .d1(q_21_26),
    .q(q_22_26)
  );
  

  flop_with_mux u_22_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_26),
    .d1(q_21_27),
    .q(q_22_27)
  );
  

  flop_with_mux u_22_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_27),
    .d1(q_21_28),
    .q(q_22_28)
  );
  

  flop_with_mux u_22_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_28),
    .d1(q_21_29),
    .q(q_22_29)
  );
  

  flop_with_mux u_22_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_29),
    .d1(q_21_30),
    .q(q_22_30)
  );
  

  flop_with_mux u_22_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_30),
    .d1(q_21_31),
    .q(q_22_31)
  );
  

  flop_with_mux u_22_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_31),
    .d1(q_21_32),
    .q(q_22_32)
  );
  

  flop_with_mux u_22_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_32),
    .d1(q_21_33),
    .q(q_22_33)
  );
  

  flop_with_mux u_22_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_33),
    .d1(q_21_34),
    .q(q_22_34)
  );
  

  flop_with_mux u_22_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_34),
    .d1(q_21_35),
    .q(q_22_35)
  );
  

  flop_with_mux u_22_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_35),
    .d1(q_21_36),
    .q(q_22_36)
  );
  

  flop_with_mux u_22_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_36),
    .d1(q_21_37),
    .q(q_22_37)
  );
  

  flop_with_mux u_22_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_37),
    .d1(q_21_38),
    .q(q_22_38)
  );
  

  flop_with_mux u_22_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_38),
    .d1(q_21_39),
    .q(q_22_39)
  );
  

  flop_with_mux u_23_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_minus1),
    .d1(q_22_0),
    .q(q_23_0)
  );
  

  flop_with_mux u_23_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_0),
    .d1(q_22_1),
    .q(q_23_1)
  );
  

  flop_with_mux u_23_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_1),
    .d1(q_22_2),
    .q(q_23_2)
  );
  

  flop_with_mux u_23_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_2),
    .d1(q_22_3),
    .q(q_23_3)
  );
  

  flop_with_mux u_23_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_3),
    .d1(q_22_4),
    .q(q_23_4)
  );
  

  flop_with_mux u_23_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_4),
    .d1(q_22_5),
    .q(q_23_5)
  );
  

  flop_with_mux u_23_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_5),
    .d1(q_22_6),
    .q(q_23_6)
  );
  

  flop_with_mux u_23_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_6),
    .d1(q_22_7),
    .q(q_23_7)
  );
  

  flop_with_mux u_23_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_7),
    .d1(q_22_8),
    .q(q_23_8)
  );
  

  flop_with_mux u_23_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_8),
    .d1(q_22_9),
    .q(q_23_9)
  );
  

  flop_with_mux u_23_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_9),
    .d1(q_22_10),
    .q(q_23_10)
  );
  

  flop_with_mux u_23_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_10),
    .d1(q_22_11),
    .q(q_23_11)
  );
  

  flop_with_mux u_23_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_11),
    .d1(q_22_12),
    .q(q_23_12)
  );
  

  flop_with_mux u_23_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_12),
    .d1(q_22_13),
    .q(q_23_13)
  );
  

  flop_with_mux u_23_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_13),
    .d1(q_22_14),
    .q(q_23_14)
  );
  

  flop_with_mux u_23_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_14),
    .d1(q_22_15),
    .q(q_23_15)
  );
  

  flop_with_mux u_23_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_15),
    .d1(q_22_16),
    .q(q_23_16)
  );
  

  flop_with_mux u_23_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_16),
    .d1(q_22_17),
    .q(q_23_17)
  );
  

  flop_with_mux u_23_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_17),
    .d1(q_22_18),
    .q(q_23_18)
  );
  

  flop_with_mux u_23_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_18),
    .d1(q_22_19),
    .q(q_23_19)
  );
  

  flop_with_mux u_23_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_19),
    .d1(q_22_20),
    .q(q_23_20)
  );
  

  flop_with_mux u_23_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_20),
    .d1(q_22_21),
    .q(q_23_21)
  );
  

  flop_with_mux u_23_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_21),
    .d1(q_22_22),
    .q(q_23_22)
  );
  

  flop_with_mux u_23_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_22),
    .d1(q_22_23),
    .q(q_23_23)
  );
  

  flop_with_mux u_23_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_23),
    .d1(q_22_24),
    .q(q_23_24)
  );
  

  flop_with_mux u_23_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_24),
    .d1(q_22_25),
    .q(q_23_25)
  );
  

  flop_with_mux u_23_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_25),
    .d1(q_22_26),
    .q(q_23_26)
  );
  

  flop_with_mux u_23_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_26),
    .d1(q_22_27),
    .q(q_23_27)
  );
  

  flop_with_mux u_23_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_27),
    .d1(q_22_28),
    .q(q_23_28)
  );
  

  flop_with_mux u_23_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_28),
    .d1(q_22_29),
    .q(q_23_29)
  );
  

  flop_with_mux u_23_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_29),
    .d1(q_22_30),
    .q(q_23_30)
  );
  

  flop_with_mux u_23_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_30),
    .d1(q_22_31),
    .q(q_23_31)
  );
  

  flop_with_mux u_23_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_31),
    .d1(q_22_32),
    .q(q_23_32)
  );
  

  flop_with_mux u_23_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_32),
    .d1(q_22_33),
    .q(q_23_33)
  );
  

  flop_with_mux u_23_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_33),
    .d1(q_22_34),
    .q(q_23_34)
  );
  

  flop_with_mux u_23_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_34),
    .d1(q_22_35),
    .q(q_23_35)
  );
  

  flop_with_mux u_23_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_35),
    .d1(q_22_36),
    .q(q_23_36)
  );
  

  flop_with_mux u_23_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_36),
    .d1(q_22_37),
    .q(q_23_37)
  );
  

  flop_with_mux u_23_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_37),
    .d1(q_22_38),
    .q(q_23_38)
  );
  

  flop_with_mux u_23_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_38),
    .d1(q_22_39),
    .q(q_23_39)
  );
  

  flop_with_mux u_24_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_minus1),
    .d1(q_23_0),
    .q(q_24_0)
  );
  

  flop_with_mux u_24_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_0),
    .d1(q_23_1),
    .q(q_24_1)
  );
  

  flop_with_mux u_24_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_1),
    .d1(q_23_2),
    .q(q_24_2)
  );
  

  flop_with_mux u_24_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_2),
    .d1(q_23_3),
    .q(q_24_3)
  );
  

  flop_with_mux u_24_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_3),
    .d1(q_23_4),
    .q(q_24_4)
  );
  

  flop_with_mux u_24_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_4),
    .d1(q_23_5),
    .q(q_24_5)
  );
  

  flop_with_mux u_24_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_5),
    .d1(q_23_6),
    .q(q_24_6)
  );
  

  flop_with_mux u_24_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_6),
    .d1(q_23_7),
    .q(q_24_7)
  );
  

  flop_with_mux u_24_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_7),
    .d1(q_23_8),
    .q(q_24_8)
  );
  

  flop_with_mux u_24_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_8),
    .d1(q_23_9),
    .q(q_24_9)
  );
  

  flop_with_mux u_24_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_9),
    .d1(q_23_10),
    .q(q_24_10)
  );
  

  flop_with_mux u_24_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_10),
    .d1(q_23_11),
    .q(q_24_11)
  );
  

  flop_with_mux u_24_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_11),
    .d1(q_23_12),
    .q(q_24_12)
  );
  

  flop_with_mux u_24_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_12),
    .d1(q_23_13),
    .q(q_24_13)
  );
  

  flop_with_mux u_24_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_13),
    .d1(q_23_14),
    .q(q_24_14)
  );
  

  flop_with_mux u_24_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_14),
    .d1(q_23_15),
    .q(q_24_15)
  );
  

  flop_with_mux u_24_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_15),
    .d1(q_23_16),
    .q(q_24_16)
  );
  

  flop_with_mux u_24_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_16),
    .d1(q_23_17),
    .q(q_24_17)
  );
  

  flop_with_mux u_24_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_17),
    .d1(q_23_18),
    .q(q_24_18)
  );
  

  flop_with_mux u_24_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_18),
    .d1(q_23_19),
    .q(q_24_19)
  );
  

  flop_with_mux u_24_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_19),
    .d1(q_23_20),
    .q(q_24_20)
  );
  

  flop_with_mux u_24_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_20),
    .d1(q_23_21),
    .q(q_24_21)
  );
  

  flop_with_mux u_24_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_21),
    .d1(q_23_22),
    .q(q_24_22)
  );
  

  flop_with_mux u_24_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_22),
    .d1(q_23_23),
    .q(q_24_23)
  );
  

  flop_with_mux u_24_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_23),
    .d1(q_23_24),
    .q(q_24_24)
  );
  

  flop_with_mux u_24_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_24),
    .d1(q_23_25),
    .q(q_24_25)
  );
  

  flop_with_mux u_24_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_25),
    .d1(q_23_26),
    .q(q_24_26)
  );
  

  flop_with_mux u_24_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_26),
    .d1(q_23_27),
    .q(q_24_27)
  );
  

  flop_with_mux u_24_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_27),
    .d1(q_23_28),
    .q(q_24_28)
  );
  

  flop_with_mux u_24_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_28),
    .d1(q_23_29),
    .q(q_24_29)
  );
  

  flop_with_mux u_24_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_29),
    .d1(q_23_30),
    .q(q_24_30)
  );
  

  flop_with_mux u_24_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_30),
    .d1(q_23_31),
    .q(q_24_31)
  );
  

  flop_with_mux u_24_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_31),
    .d1(q_23_32),
    .q(q_24_32)
  );
  

  flop_with_mux u_24_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_32),
    .d1(q_23_33),
    .q(q_24_33)
  );
  

  flop_with_mux u_24_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_33),
    .d1(q_23_34),
    .q(q_24_34)
  );
  

  flop_with_mux u_24_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_34),
    .d1(q_23_35),
    .q(q_24_35)
  );
  

  flop_with_mux u_24_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_35),
    .d1(q_23_36),
    .q(q_24_36)
  );
  

  flop_with_mux u_24_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_36),
    .d1(q_23_37),
    .q(q_24_37)
  );
  

  flop_with_mux u_24_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_37),
    .d1(q_23_38),
    .q(q_24_38)
  );
  

  flop_with_mux u_24_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_38),
    .d1(q_23_39),
    .q(q_24_39)
  );
  

  flop_with_mux u_25_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_minus1),
    .d1(q_24_0),
    .q(q_25_0)
  );
  

  flop_with_mux u_25_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_0),
    .d1(q_24_1),
    .q(q_25_1)
  );
  

  flop_with_mux u_25_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_1),
    .d1(q_24_2),
    .q(q_25_2)
  );
  

  flop_with_mux u_25_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_2),
    .d1(q_24_3),
    .q(q_25_3)
  );
  

  flop_with_mux u_25_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_3),
    .d1(q_24_4),
    .q(q_25_4)
  );
  

  flop_with_mux u_25_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_4),
    .d1(q_24_5),
    .q(q_25_5)
  );
  

  flop_with_mux u_25_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_5),
    .d1(q_24_6),
    .q(q_25_6)
  );
  

  flop_with_mux u_25_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_6),
    .d1(q_24_7),
    .q(q_25_7)
  );
  

  flop_with_mux u_25_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_7),
    .d1(q_24_8),
    .q(q_25_8)
  );
  

  flop_with_mux u_25_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_8),
    .d1(q_24_9),
    .q(q_25_9)
  );
  

  flop_with_mux u_25_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_9),
    .d1(q_24_10),
    .q(q_25_10)
  );
  

  flop_with_mux u_25_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_10),
    .d1(q_24_11),
    .q(q_25_11)
  );
  

  flop_with_mux u_25_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_11),
    .d1(q_24_12),
    .q(q_25_12)
  );
  

  flop_with_mux u_25_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_12),
    .d1(q_24_13),
    .q(q_25_13)
  );
  

  flop_with_mux u_25_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_13),
    .d1(q_24_14),
    .q(q_25_14)
  );
  

  flop_with_mux u_25_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_14),
    .d1(q_24_15),
    .q(q_25_15)
  );
  

  flop_with_mux u_25_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_15),
    .d1(q_24_16),
    .q(q_25_16)
  );
  

  flop_with_mux u_25_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_16),
    .d1(q_24_17),
    .q(q_25_17)
  );
  

  flop_with_mux u_25_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_17),
    .d1(q_24_18),
    .q(q_25_18)
  );
  

  flop_with_mux u_25_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_18),
    .d1(q_24_19),
    .q(q_25_19)
  );
  

  flop_with_mux u_25_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_19),
    .d1(q_24_20),
    .q(q_25_20)
  );
  

  flop_with_mux u_25_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_20),
    .d1(q_24_21),
    .q(q_25_21)
  );
  

  flop_with_mux u_25_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_21),
    .d1(q_24_22),
    .q(q_25_22)
  );
  

  flop_with_mux u_25_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_22),
    .d1(q_24_23),
    .q(q_25_23)
  );
  

  flop_with_mux u_25_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_23),
    .d1(q_24_24),
    .q(q_25_24)
  );
  

  flop_with_mux u_25_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_24),
    .d1(q_24_25),
    .q(q_25_25)
  );
  

  flop_with_mux u_25_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_25),
    .d1(q_24_26),
    .q(q_25_26)
  );
  

  flop_with_mux u_25_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_26),
    .d1(q_24_27),
    .q(q_25_27)
  );
  

  flop_with_mux u_25_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_27),
    .d1(q_24_28),
    .q(q_25_28)
  );
  

  flop_with_mux u_25_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_28),
    .d1(q_24_29),
    .q(q_25_29)
  );
  

  flop_with_mux u_25_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_29),
    .d1(q_24_30),
    .q(q_25_30)
  );
  

  flop_with_mux u_25_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_30),
    .d1(q_24_31),
    .q(q_25_31)
  );
  

  flop_with_mux u_25_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_31),
    .d1(q_24_32),
    .q(q_25_32)
  );
  

  flop_with_mux u_25_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_32),
    .d1(q_24_33),
    .q(q_25_33)
  );
  

  flop_with_mux u_25_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_33),
    .d1(q_24_34),
    .q(q_25_34)
  );
  

  flop_with_mux u_25_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_34),
    .d1(q_24_35),
    .q(q_25_35)
  );
  

  flop_with_mux u_25_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_35),
    .d1(q_24_36),
    .q(q_25_36)
  );
  

  flop_with_mux u_25_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_36),
    .d1(q_24_37),
    .q(q_25_37)
  );
  

  flop_with_mux u_25_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_37),
    .d1(q_24_38),
    .q(q_25_38)
  );
  

  flop_with_mux u_25_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_38),
    .d1(q_24_39),
    .q(q_25_39)
  );
  

  flop_with_mux u_26_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_minus1),
    .d1(q_25_0),
    .q(q_26_0)
  );
  

  flop_with_mux u_26_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_0),
    .d1(q_25_1),
    .q(q_26_1)
  );
  

  flop_with_mux u_26_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_1),
    .d1(q_25_2),
    .q(q_26_2)
  );
  

  flop_with_mux u_26_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_2),
    .d1(q_25_3),
    .q(q_26_3)
  );
  

  flop_with_mux u_26_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_3),
    .d1(q_25_4),
    .q(q_26_4)
  );
  

  flop_with_mux u_26_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_4),
    .d1(q_25_5),
    .q(q_26_5)
  );
  

  flop_with_mux u_26_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_5),
    .d1(q_25_6),
    .q(q_26_6)
  );
  

  flop_with_mux u_26_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_6),
    .d1(q_25_7),
    .q(q_26_7)
  );
  

  flop_with_mux u_26_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_7),
    .d1(q_25_8),
    .q(q_26_8)
  );
  

  flop_with_mux u_26_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_8),
    .d1(q_25_9),
    .q(q_26_9)
  );
  

  flop_with_mux u_26_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_9),
    .d1(q_25_10),
    .q(q_26_10)
  );
  

  flop_with_mux u_26_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_10),
    .d1(q_25_11),
    .q(q_26_11)
  );
  

  flop_with_mux u_26_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_11),
    .d1(q_25_12),
    .q(q_26_12)
  );
  

  flop_with_mux u_26_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_12),
    .d1(q_25_13),
    .q(q_26_13)
  );
  

  flop_with_mux u_26_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_13),
    .d1(q_25_14),
    .q(q_26_14)
  );
  

  flop_with_mux u_26_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_14),
    .d1(q_25_15),
    .q(q_26_15)
  );
  

  flop_with_mux u_26_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_15),
    .d1(q_25_16),
    .q(q_26_16)
  );
  

  flop_with_mux u_26_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_16),
    .d1(q_25_17),
    .q(q_26_17)
  );
  

  flop_with_mux u_26_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_17),
    .d1(q_25_18),
    .q(q_26_18)
  );
  

  flop_with_mux u_26_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_18),
    .d1(q_25_19),
    .q(q_26_19)
  );
  

  flop_with_mux u_26_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_19),
    .d1(q_25_20),
    .q(q_26_20)
  );
  

  flop_with_mux u_26_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_20),
    .d1(q_25_21),
    .q(q_26_21)
  );
  

  flop_with_mux u_26_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_21),
    .d1(q_25_22),
    .q(q_26_22)
  );
  

  flop_with_mux u_26_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_22),
    .d1(q_25_23),
    .q(q_26_23)
  );
  

  flop_with_mux u_26_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_23),
    .d1(q_25_24),
    .q(q_26_24)
  );
  

  flop_with_mux u_26_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_24),
    .d1(q_25_25),
    .q(q_26_25)
  );
  

  flop_with_mux u_26_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_25),
    .d1(q_25_26),
    .q(q_26_26)
  );
  

  flop_with_mux u_26_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_26),
    .d1(q_25_27),
    .q(q_26_27)
  );
  

  flop_with_mux u_26_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_27),
    .d1(q_25_28),
    .q(q_26_28)
  );
  

  flop_with_mux u_26_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_28),
    .d1(q_25_29),
    .q(q_26_29)
  );
  

  flop_with_mux u_26_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_29),
    .d1(q_25_30),
    .q(q_26_30)
  );
  

  flop_with_mux u_26_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_30),
    .d1(q_25_31),
    .q(q_26_31)
  );
  

  flop_with_mux u_26_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_31),
    .d1(q_25_32),
    .q(q_26_32)
  );
  

  flop_with_mux u_26_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_32),
    .d1(q_25_33),
    .q(q_26_33)
  );
  

  flop_with_mux u_26_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_33),
    .d1(q_25_34),
    .q(q_26_34)
  );
  

  flop_with_mux u_26_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_34),
    .d1(q_25_35),
    .q(q_26_35)
  );
  

  flop_with_mux u_26_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_35),
    .d1(q_25_36),
    .q(q_26_36)
  );
  

  flop_with_mux u_26_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_36),
    .d1(q_25_37),
    .q(q_26_37)
  );
  

  flop_with_mux u_26_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_37),
    .d1(q_25_38),
    .q(q_26_38)
  );
  

  flop_with_mux u_26_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_38),
    .d1(q_25_39),
    .q(q_26_39)
  );
  

  flop_with_mux u_27_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_minus1),
    .d1(q_26_0),
    .q(q_27_0)
  );
  

  flop_with_mux u_27_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_0),
    .d1(q_26_1),
    .q(q_27_1)
  );
  

  flop_with_mux u_27_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_1),
    .d1(q_26_2),
    .q(q_27_2)
  );
  

  flop_with_mux u_27_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_2),
    .d1(q_26_3),
    .q(q_27_3)
  );
  

  flop_with_mux u_27_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_3),
    .d1(q_26_4),
    .q(q_27_4)
  );
  

  flop_with_mux u_27_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_4),
    .d1(q_26_5),
    .q(q_27_5)
  );
  

  flop_with_mux u_27_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_5),
    .d1(q_26_6),
    .q(q_27_6)
  );
  

  flop_with_mux u_27_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_6),
    .d1(q_26_7),
    .q(q_27_7)
  );
  

  flop_with_mux u_27_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_7),
    .d1(q_26_8),
    .q(q_27_8)
  );
  

  flop_with_mux u_27_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_8),
    .d1(q_26_9),
    .q(q_27_9)
  );
  

  flop_with_mux u_27_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_9),
    .d1(q_26_10),
    .q(q_27_10)
  );
  

  flop_with_mux u_27_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_10),
    .d1(q_26_11),
    .q(q_27_11)
  );
  

  flop_with_mux u_27_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_11),
    .d1(q_26_12),
    .q(q_27_12)
  );
  

  flop_with_mux u_27_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_12),
    .d1(q_26_13),
    .q(q_27_13)
  );
  

  flop_with_mux u_27_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_13),
    .d1(q_26_14),
    .q(q_27_14)
  );
  

  flop_with_mux u_27_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_14),
    .d1(q_26_15),
    .q(q_27_15)
  );
  

  flop_with_mux u_27_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_15),
    .d1(q_26_16),
    .q(q_27_16)
  );
  

  flop_with_mux u_27_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_16),
    .d1(q_26_17),
    .q(q_27_17)
  );
  

  flop_with_mux u_27_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_17),
    .d1(q_26_18),
    .q(q_27_18)
  );
  

  flop_with_mux u_27_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_18),
    .d1(q_26_19),
    .q(q_27_19)
  );
  

  flop_with_mux u_27_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_19),
    .d1(q_26_20),
    .q(q_27_20)
  );
  

  flop_with_mux u_27_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_20),
    .d1(q_26_21),
    .q(q_27_21)
  );
  

  flop_with_mux u_27_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_21),
    .d1(q_26_22),
    .q(q_27_22)
  );
  

  flop_with_mux u_27_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_22),
    .d1(q_26_23),
    .q(q_27_23)
  );
  

  flop_with_mux u_27_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_23),
    .d1(q_26_24),
    .q(q_27_24)
  );
  

  flop_with_mux u_27_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_24),
    .d1(q_26_25),
    .q(q_27_25)
  );
  

  flop_with_mux u_27_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_25),
    .d1(q_26_26),
    .q(q_27_26)
  );
  

  flop_with_mux u_27_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_26),
    .d1(q_26_27),
    .q(q_27_27)
  );
  

  flop_with_mux u_27_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_27),
    .d1(q_26_28),
    .q(q_27_28)
  );
  

  flop_with_mux u_27_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_28),
    .d1(q_26_29),
    .q(q_27_29)
  );
  

  flop_with_mux u_27_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_29),
    .d1(q_26_30),
    .q(q_27_30)
  );
  

  flop_with_mux u_27_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_30),
    .d1(q_26_31),
    .q(q_27_31)
  );
  

  flop_with_mux u_27_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_31),
    .d1(q_26_32),
    .q(q_27_32)
  );
  

  flop_with_mux u_27_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_32),
    .d1(q_26_33),
    .q(q_27_33)
  );
  

  flop_with_mux u_27_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_33),
    .d1(q_26_34),
    .q(q_27_34)
  );
  

  flop_with_mux u_27_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_34),
    .d1(q_26_35),
    .q(q_27_35)
  );
  

  flop_with_mux u_27_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_35),
    .d1(q_26_36),
    .q(q_27_36)
  );
  

  flop_with_mux u_27_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_36),
    .d1(q_26_37),
    .q(q_27_37)
  );
  

  flop_with_mux u_27_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_37),
    .d1(q_26_38),
    .q(q_27_38)
  );
  

  flop_with_mux u_27_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_38),
    .d1(q_26_39),
    .q(q_27_39)
  );
  

  flop_with_mux u_28_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_minus1),
    .d1(q_27_0),
    .q(q_28_0)
  );
  

  flop_with_mux u_28_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_0),
    .d1(q_27_1),
    .q(q_28_1)
  );
  

  flop_with_mux u_28_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_1),
    .d1(q_27_2),
    .q(q_28_2)
  );
  

  flop_with_mux u_28_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_2),
    .d1(q_27_3),
    .q(q_28_3)
  );
  

  flop_with_mux u_28_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_3),
    .d1(q_27_4),
    .q(q_28_4)
  );
  

  flop_with_mux u_28_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_4),
    .d1(q_27_5),
    .q(q_28_5)
  );
  

  flop_with_mux u_28_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_5),
    .d1(q_27_6),
    .q(q_28_6)
  );
  

  flop_with_mux u_28_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_6),
    .d1(q_27_7),
    .q(q_28_7)
  );
  

  flop_with_mux u_28_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_7),
    .d1(q_27_8),
    .q(q_28_8)
  );
  

  flop_with_mux u_28_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_8),
    .d1(q_27_9),
    .q(q_28_9)
  );
  

  flop_with_mux u_28_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_9),
    .d1(q_27_10),
    .q(q_28_10)
  );
  

  flop_with_mux u_28_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_10),
    .d1(q_27_11),
    .q(q_28_11)
  );
  

  flop_with_mux u_28_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_11),
    .d1(q_27_12),
    .q(q_28_12)
  );
  

  flop_with_mux u_28_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_12),
    .d1(q_27_13),
    .q(q_28_13)
  );
  

  flop_with_mux u_28_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_13),
    .d1(q_27_14),
    .q(q_28_14)
  );
  

  flop_with_mux u_28_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_14),
    .d1(q_27_15),
    .q(q_28_15)
  );
  

  flop_with_mux u_28_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_15),
    .d1(q_27_16),
    .q(q_28_16)
  );
  

  flop_with_mux u_28_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_16),
    .d1(q_27_17),
    .q(q_28_17)
  );
  

  flop_with_mux u_28_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_17),
    .d1(q_27_18),
    .q(q_28_18)
  );
  

  flop_with_mux u_28_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_18),
    .d1(q_27_19),
    .q(q_28_19)
  );
  

  flop_with_mux u_28_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_19),
    .d1(q_27_20),
    .q(q_28_20)
  );
  

  flop_with_mux u_28_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_20),
    .d1(q_27_21),
    .q(q_28_21)
  );
  

  flop_with_mux u_28_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_21),
    .d1(q_27_22),
    .q(q_28_22)
  );
  

  flop_with_mux u_28_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_22),
    .d1(q_27_23),
    .q(q_28_23)
  );
  

  flop_with_mux u_28_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_23),
    .d1(q_27_24),
    .q(q_28_24)
  );
  

  flop_with_mux u_28_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_24),
    .d1(q_27_25),
    .q(q_28_25)
  );
  

  flop_with_mux u_28_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_25),
    .d1(q_27_26),
    .q(q_28_26)
  );
  

  flop_with_mux u_28_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_26),
    .d1(q_27_27),
    .q(q_28_27)
  );
  

  flop_with_mux u_28_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_27),
    .d1(q_27_28),
    .q(q_28_28)
  );
  

  flop_with_mux u_28_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_28),
    .d1(q_27_29),
    .q(q_28_29)
  );
  

  flop_with_mux u_28_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_29),
    .d1(q_27_30),
    .q(q_28_30)
  );
  

  flop_with_mux u_28_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_30),
    .d1(q_27_31),
    .q(q_28_31)
  );
  

  flop_with_mux u_28_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_31),
    .d1(q_27_32),
    .q(q_28_32)
  );
  

  flop_with_mux u_28_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_32),
    .d1(q_27_33),
    .q(q_28_33)
  );
  

  flop_with_mux u_28_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_33),
    .d1(q_27_34),
    .q(q_28_34)
  );
  

  flop_with_mux u_28_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_34),
    .d1(q_27_35),
    .q(q_28_35)
  );
  

  flop_with_mux u_28_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_35),
    .d1(q_27_36),
    .q(q_28_36)
  );
  

  flop_with_mux u_28_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_36),
    .d1(q_27_37),
    .q(q_28_37)
  );
  

  flop_with_mux u_28_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_37),
    .d1(q_27_38),
    .q(q_28_38)
  );
  

  flop_with_mux u_28_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_38),
    .d1(q_27_39),
    .q(q_28_39)
  );
  

  flop_with_mux u_29_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_minus1),
    .d1(q_28_0),
    .q(q_29_0)
  );
  

  flop_with_mux u_29_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_0),
    .d1(q_28_1),
    .q(q_29_1)
  );
  

  flop_with_mux u_29_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_1),
    .d1(q_28_2),
    .q(q_29_2)
  );
  

  flop_with_mux u_29_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_2),
    .d1(q_28_3),
    .q(q_29_3)
  );
  

  flop_with_mux u_29_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_3),
    .d1(q_28_4),
    .q(q_29_4)
  );
  

  flop_with_mux u_29_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_4),
    .d1(q_28_5),
    .q(q_29_5)
  );
  

  flop_with_mux u_29_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_5),
    .d1(q_28_6),
    .q(q_29_6)
  );
  

  flop_with_mux u_29_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_6),
    .d1(q_28_7),
    .q(q_29_7)
  );
  

  flop_with_mux u_29_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_7),
    .d1(q_28_8),
    .q(q_29_8)
  );
  

  flop_with_mux u_29_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_8),
    .d1(q_28_9),
    .q(q_29_9)
  );
  

  flop_with_mux u_29_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_9),
    .d1(q_28_10),
    .q(q_29_10)
  );
  

  flop_with_mux u_29_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_10),
    .d1(q_28_11),
    .q(q_29_11)
  );
  

  flop_with_mux u_29_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_11),
    .d1(q_28_12),
    .q(q_29_12)
  );
  

  flop_with_mux u_29_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_12),
    .d1(q_28_13),
    .q(q_29_13)
  );
  

  flop_with_mux u_29_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_13),
    .d1(q_28_14),
    .q(q_29_14)
  );
  

  flop_with_mux u_29_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_14),
    .d1(q_28_15),
    .q(q_29_15)
  );
  

  flop_with_mux u_29_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_15),
    .d1(q_28_16),
    .q(q_29_16)
  );
  

  flop_with_mux u_29_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_16),
    .d1(q_28_17),
    .q(q_29_17)
  );
  

  flop_with_mux u_29_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_17),
    .d1(q_28_18),
    .q(q_29_18)
  );
  

  flop_with_mux u_29_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_18),
    .d1(q_28_19),
    .q(q_29_19)
  );
  

  flop_with_mux u_29_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_19),
    .d1(q_28_20),
    .q(q_29_20)
  );
  

  flop_with_mux u_29_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_20),
    .d1(q_28_21),
    .q(q_29_21)
  );
  

  flop_with_mux u_29_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_21),
    .d1(q_28_22),
    .q(q_29_22)
  );
  

  flop_with_mux u_29_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_22),
    .d1(q_28_23),
    .q(q_29_23)
  );
  

  flop_with_mux u_29_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_23),
    .d1(q_28_24),
    .q(q_29_24)
  );
  

  flop_with_mux u_29_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_24),
    .d1(q_28_25),
    .q(q_29_25)
  );
  

  flop_with_mux u_29_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_25),
    .d1(q_28_26),
    .q(q_29_26)
  );
  

  flop_with_mux u_29_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_26),
    .d1(q_28_27),
    .q(q_29_27)
  );
  

  flop_with_mux u_29_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_27),
    .d1(q_28_28),
    .q(q_29_28)
  );
  

  flop_with_mux u_29_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_28),
    .d1(q_28_29),
    .q(q_29_29)
  );
  

  flop_with_mux u_29_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_29),
    .d1(q_28_30),
    .q(q_29_30)
  );
  

  flop_with_mux u_29_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_30),
    .d1(q_28_31),
    .q(q_29_31)
  );
  

  flop_with_mux u_29_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_31),
    .d1(q_28_32),
    .q(q_29_32)
  );
  

  flop_with_mux u_29_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_32),
    .d1(q_28_33),
    .q(q_29_33)
  );
  

  flop_with_mux u_29_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_33),
    .d1(q_28_34),
    .q(q_29_34)
  );
  

  flop_with_mux u_29_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_34),
    .d1(q_28_35),
    .q(q_29_35)
  );
  

  flop_with_mux u_29_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_35),
    .d1(q_28_36),
    .q(q_29_36)
  );
  

  flop_with_mux u_29_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_36),
    .d1(q_28_37),
    .q(q_29_37)
  );
  

  flop_with_mux u_29_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_37),
    .d1(q_28_38),
    .q(q_29_38)
  );
  

  flop_with_mux u_29_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_38),
    .d1(q_28_39),
    .q(q_29_39)
  );
  

  flop_with_mux u_30_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_minus1),
    .d1(q_29_0),
    .q(q_30_0)
  );
  

  flop_with_mux u_30_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_0),
    .d1(q_29_1),
    .q(q_30_1)
  );
  

  flop_with_mux u_30_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_1),
    .d1(q_29_2),
    .q(q_30_2)
  );
  

  flop_with_mux u_30_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_2),
    .d1(q_29_3),
    .q(q_30_3)
  );
  

  flop_with_mux u_30_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_3),
    .d1(q_29_4),
    .q(q_30_4)
  );
  

  flop_with_mux u_30_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_4),
    .d1(q_29_5),
    .q(q_30_5)
  );
  

  flop_with_mux u_30_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_5),
    .d1(q_29_6),
    .q(q_30_6)
  );
  

  flop_with_mux u_30_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_6),
    .d1(q_29_7),
    .q(q_30_7)
  );
  

  flop_with_mux u_30_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_7),
    .d1(q_29_8),
    .q(q_30_8)
  );
  

  flop_with_mux u_30_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_8),
    .d1(q_29_9),
    .q(q_30_9)
  );
  

  flop_with_mux u_30_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_9),
    .d1(q_29_10),
    .q(q_30_10)
  );
  

  flop_with_mux u_30_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_10),
    .d1(q_29_11),
    .q(q_30_11)
  );
  

  flop_with_mux u_30_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_11),
    .d1(q_29_12),
    .q(q_30_12)
  );
  

  flop_with_mux u_30_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_12),
    .d1(q_29_13),
    .q(q_30_13)
  );
  

  flop_with_mux u_30_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_13),
    .d1(q_29_14),
    .q(q_30_14)
  );
  

  flop_with_mux u_30_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_14),
    .d1(q_29_15),
    .q(q_30_15)
  );
  

  flop_with_mux u_30_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_15),
    .d1(q_29_16),
    .q(q_30_16)
  );
  

  flop_with_mux u_30_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_16),
    .d1(q_29_17),
    .q(q_30_17)
  );
  

  flop_with_mux u_30_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_17),
    .d1(q_29_18),
    .q(q_30_18)
  );
  

  flop_with_mux u_30_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_18),
    .d1(q_29_19),
    .q(q_30_19)
  );
  

  flop_with_mux u_30_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_19),
    .d1(q_29_20),
    .q(q_30_20)
  );
  

  flop_with_mux u_30_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_20),
    .d1(q_29_21),
    .q(q_30_21)
  );
  

  flop_with_mux u_30_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_21),
    .d1(q_29_22),
    .q(q_30_22)
  );
  

  flop_with_mux u_30_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_22),
    .d1(q_29_23),
    .q(q_30_23)
  );
  

  flop_with_mux u_30_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_23),
    .d1(q_29_24),
    .q(q_30_24)
  );
  

  flop_with_mux u_30_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_24),
    .d1(q_29_25),
    .q(q_30_25)
  );
  

  flop_with_mux u_30_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_25),
    .d1(q_29_26),
    .q(q_30_26)
  );
  

  flop_with_mux u_30_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_26),
    .d1(q_29_27),
    .q(q_30_27)
  );
  

  flop_with_mux u_30_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_27),
    .d1(q_29_28),
    .q(q_30_28)
  );
  

  flop_with_mux u_30_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_28),
    .d1(q_29_29),
    .q(q_30_29)
  );
  

  flop_with_mux u_30_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_29),
    .d1(q_29_30),
    .q(q_30_30)
  );
  

  flop_with_mux u_30_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_30),
    .d1(q_29_31),
    .q(q_30_31)
  );
  

  flop_with_mux u_30_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_31),
    .d1(q_29_32),
    .q(q_30_32)
  );
  

  flop_with_mux u_30_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_32),
    .d1(q_29_33),
    .q(q_30_33)
  );
  

  flop_with_mux u_30_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_33),
    .d1(q_29_34),
    .q(q_30_34)
  );
  

  flop_with_mux u_30_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_34),
    .d1(q_29_35),
    .q(q_30_35)
  );
  

  flop_with_mux u_30_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_35),
    .d1(q_29_36),
    .q(q_30_36)
  );
  

  flop_with_mux u_30_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_36),
    .d1(q_29_37),
    .q(q_30_37)
  );
  

  flop_with_mux u_30_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_37),
    .d1(q_29_38),
    .q(q_30_38)
  );
  

  flop_with_mux u_30_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_38),
    .d1(q_29_39),
    .q(q_30_39)
  );
  

  flop_with_mux u_31_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_minus1),
    .d1(q_30_0),
    .q(q_31_0)
  );
  

  flop_with_mux u_31_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_0),
    .d1(q_30_1),
    .q(q_31_1)
  );
  

  flop_with_mux u_31_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_1),
    .d1(q_30_2),
    .q(q_31_2)
  );
  

  flop_with_mux u_31_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_2),
    .d1(q_30_3),
    .q(q_31_3)
  );
  

  flop_with_mux u_31_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_3),
    .d1(q_30_4),
    .q(q_31_4)
  );
  

  flop_with_mux u_31_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_4),
    .d1(q_30_5),
    .q(q_31_5)
  );
  

  flop_with_mux u_31_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_5),
    .d1(q_30_6),
    .q(q_31_6)
  );
  

  flop_with_mux u_31_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_6),
    .d1(q_30_7),
    .q(q_31_7)
  );
  

  flop_with_mux u_31_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_7),
    .d1(q_30_8),
    .q(q_31_8)
  );
  

  flop_with_mux u_31_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_8),
    .d1(q_30_9),
    .q(q_31_9)
  );
  

  flop_with_mux u_31_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_9),
    .d1(q_30_10),
    .q(q_31_10)
  );
  

  flop_with_mux u_31_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_10),
    .d1(q_30_11),
    .q(q_31_11)
  );
  

  flop_with_mux u_31_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_11),
    .d1(q_30_12),
    .q(q_31_12)
  );
  

  flop_with_mux u_31_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_12),
    .d1(q_30_13),
    .q(q_31_13)
  );
  

  flop_with_mux u_31_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_13),
    .d1(q_30_14),
    .q(q_31_14)
  );
  

  flop_with_mux u_31_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_14),
    .d1(q_30_15),
    .q(q_31_15)
  );
  

  flop_with_mux u_31_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_15),
    .d1(q_30_16),
    .q(q_31_16)
  );
  

  flop_with_mux u_31_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_16),
    .d1(q_30_17),
    .q(q_31_17)
  );
  

  flop_with_mux u_31_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_17),
    .d1(q_30_18),
    .q(q_31_18)
  );
  

  flop_with_mux u_31_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_18),
    .d1(q_30_19),
    .q(q_31_19)
  );
  

  flop_with_mux u_31_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_19),
    .d1(q_30_20),
    .q(q_31_20)
  );
  

  flop_with_mux u_31_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_20),
    .d1(q_30_21),
    .q(q_31_21)
  );
  

  flop_with_mux u_31_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_21),
    .d1(q_30_22),
    .q(q_31_22)
  );
  

  flop_with_mux u_31_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_22),
    .d1(q_30_23),
    .q(q_31_23)
  );
  

  flop_with_mux u_31_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_23),
    .d1(q_30_24),
    .q(q_31_24)
  );
  

  flop_with_mux u_31_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_24),
    .d1(q_30_25),
    .q(q_31_25)
  );
  

  flop_with_mux u_31_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_25),
    .d1(q_30_26),
    .q(q_31_26)
  );
  

  flop_with_mux u_31_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_26),
    .d1(q_30_27),
    .q(q_31_27)
  );
  

  flop_with_mux u_31_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_27),
    .d1(q_30_28),
    .q(q_31_28)
  );
  

  flop_with_mux u_31_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_28),
    .d1(q_30_29),
    .q(q_31_29)
  );
  

  flop_with_mux u_31_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_29),
    .d1(q_30_30),
    .q(q_31_30)
  );
  

  flop_with_mux u_31_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_30),
    .d1(q_30_31),
    .q(q_31_31)
  );
  

  flop_with_mux u_31_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_31),
    .d1(q_30_32),
    .q(q_31_32)
  );
  

  flop_with_mux u_31_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_32),
    .d1(q_30_33),
    .q(q_31_33)
  );
  

  flop_with_mux u_31_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_33),
    .d1(q_30_34),
    .q(q_31_34)
  );
  

  flop_with_mux u_31_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_34),
    .d1(q_30_35),
    .q(q_31_35)
  );
  

  flop_with_mux u_31_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_35),
    .d1(q_30_36),
    .q(q_31_36)
  );
  

  flop_with_mux u_31_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_36),
    .d1(q_30_37),
    .q(q_31_37)
  );
  

  flop_with_mux u_31_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_37),
    .d1(q_30_38),
    .q(q_31_38)
  );
  

  flop_with_mux u_31_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_38),
    .d1(q_30_39),
    .q(q_31_39)
  );
  

  flop_with_mux u_32_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_minus1),
    .d1(q_31_0),
    .q(q_32_0)
  );
  

  flop_with_mux u_32_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_0),
    .d1(q_31_1),
    .q(q_32_1)
  );
  

  flop_with_mux u_32_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_1),
    .d1(q_31_2),
    .q(q_32_2)
  );
  

  flop_with_mux u_32_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_2),
    .d1(q_31_3),
    .q(q_32_3)
  );
  

  flop_with_mux u_32_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_3),
    .d1(q_31_4),
    .q(q_32_4)
  );
  

  flop_with_mux u_32_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_4),
    .d1(q_31_5),
    .q(q_32_5)
  );
  

  flop_with_mux u_32_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_5),
    .d1(q_31_6),
    .q(q_32_6)
  );
  

  flop_with_mux u_32_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_6),
    .d1(q_31_7),
    .q(q_32_7)
  );
  

  flop_with_mux u_32_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_7),
    .d1(q_31_8),
    .q(q_32_8)
  );
  

  flop_with_mux u_32_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_8),
    .d1(q_31_9),
    .q(q_32_9)
  );
  

  flop_with_mux u_32_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_9),
    .d1(q_31_10),
    .q(q_32_10)
  );
  

  flop_with_mux u_32_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_10),
    .d1(q_31_11),
    .q(q_32_11)
  );
  

  flop_with_mux u_32_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_11),
    .d1(q_31_12),
    .q(q_32_12)
  );
  

  flop_with_mux u_32_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_12),
    .d1(q_31_13),
    .q(q_32_13)
  );
  

  flop_with_mux u_32_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_13),
    .d1(q_31_14),
    .q(q_32_14)
  );
  

  flop_with_mux u_32_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_14),
    .d1(q_31_15),
    .q(q_32_15)
  );
  

  flop_with_mux u_32_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_15),
    .d1(q_31_16),
    .q(q_32_16)
  );
  

  flop_with_mux u_32_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_16),
    .d1(q_31_17),
    .q(q_32_17)
  );
  

  flop_with_mux u_32_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_17),
    .d1(q_31_18),
    .q(q_32_18)
  );
  

  flop_with_mux u_32_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_18),
    .d1(q_31_19),
    .q(q_32_19)
  );
  

  flop_with_mux u_32_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_19),
    .d1(q_31_20),
    .q(q_32_20)
  );
  

  flop_with_mux u_32_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_20),
    .d1(q_31_21),
    .q(q_32_21)
  );
  

  flop_with_mux u_32_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_21),
    .d1(q_31_22),
    .q(q_32_22)
  );
  

  flop_with_mux u_32_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_22),
    .d1(q_31_23),
    .q(q_32_23)
  );
  

  flop_with_mux u_32_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_23),
    .d1(q_31_24),
    .q(q_32_24)
  );
  

  flop_with_mux u_32_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_24),
    .d1(q_31_25),
    .q(q_32_25)
  );
  

  flop_with_mux u_32_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_25),
    .d1(q_31_26),
    .q(q_32_26)
  );
  

  flop_with_mux u_32_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_26),
    .d1(q_31_27),
    .q(q_32_27)
  );
  

  flop_with_mux u_32_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_27),
    .d1(q_31_28),
    .q(q_32_28)
  );
  

  flop_with_mux u_32_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_28),
    .d1(q_31_29),
    .q(q_32_29)
  );
  

  flop_with_mux u_32_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_29),
    .d1(q_31_30),
    .q(q_32_30)
  );
  

  flop_with_mux u_32_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_30),
    .d1(q_31_31),
    .q(q_32_31)
  );
  

  flop_with_mux u_32_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_31),
    .d1(q_31_32),
    .q(q_32_32)
  );
  

  flop_with_mux u_32_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_32),
    .d1(q_31_33),
    .q(q_32_33)
  );
  

  flop_with_mux u_32_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_33),
    .d1(q_31_34),
    .q(q_32_34)
  );
  

  flop_with_mux u_32_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_34),
    .d1(q_31_35),
    .q(q_32_35)
  );
  

  flop_with_mux u_32_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_35),
    .d1(q_31_36),
    .q(q_32_36)
  );
  

  flop_with_mux u_32_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_36),
    .d1(q_31_37),
    .q(q_32_37)
  );
  

  flop_with_mux u_32_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_37),
    .d1(q_31_38),
    .q(q_32_38)
  );
  

  flop_with_mux u_32_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_38),
    .d1(q_31_39),
    .q(q_32_39)
  );
  

  flop_with_mux u_33_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_minus1),
    .d1(q_32_0),
    .q(q_33_0)
  );
  

  flop_with_mux u_33_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_0),
    .d1(q_32_1),
    .q(q_33_1)
  );
  

  flop_with_mux u_33_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_1),
    .d1(q_32_2),
    .q(q_33_2)
  );
  

  flop_with_mux u_33_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_2),
    .d1(q_32_3),
    .q(q_33_3)
  );
  

  flop_with_mux u_33_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_3),
    .d1(q_32_4),
    .q(q_33_4)
  );
  

  flop_with_mux u_33_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_4),
    .d1(q_32_5),
    .q(q_33_5)
  );
  

  flop_with_mux u_33_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_5),
    .d1(q_32_6),
    .q(q_33_6)
  );
  

  flop_with_mux u_33_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_6),
    .d1(q_32_7),
    .q(q_33_7)
  );
  

  flop_with_mux u_33_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_7),
    .d1(q_32_8),
    .q(q_33_8)
  );
  

  flop_with_mux u_33_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_8),
    .d1(q_32_9),
    .q(q_33_9)
  );
  

  flop_with_mux u_33_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_9),
    .d1(q_32_10),
    .q(q_33_10)
  );
  

  flop_with_mux u_33_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_10),
    .d1(q_32_11),
    .q(q_33_11)
  );
  

  flop_with_mux u_33_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_11),
    .d1(q_32_12),
    .q(q_33_12)
  );
  

  flop_with_mux u_33_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_12),
    .d1(q_32_13),
    .q(q_33_13)
  );
  

  flop_with_mux u_33_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_13),
    .d1(q_32_14),
    .q(q_33_14)
  );
  

  flop_with_mux u_33_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_14),
    .d1(q_32_15),
    .q(q_33_15)
  );
  

  flop_with_mux u_33_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_15),
    .d1(q_32_16),
    .q(q_33_16)
  );
  

  flop_with_mux u_33_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_16),
    .d1(q_32_17),
    .q(q_33_17)
  );
  

  flop_with_mux u_33_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_17),
    .d1(q_32_18),
    .q(q_33_18)
  );
  

  flop_with_mux u_33_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_18),
    .d1(q_32_19),
    .q(q_33_19)
  );
  

  flop_with_mux u_33_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_19),
    .d1(q_32_20),
    .q(q_33_20)
  );
  

  flop_with_mux u_33_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_20),
    .d1(q_32_21),
    .q(q_33_21)
  );
  

  flop_with_mux u_33_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_21),
    .d1(q_32_22),
    .q(q_33_22)
  );
  

  flop_with_mux u_33_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_22),
    .d1(q_32_23),
    .q(q_33_23)
  );
  

  flop_with_mux u_33_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_23),
    .d1(q_32_24),
    .q(q_33_24)
  );
  

  flop_with_mux u_33_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_24),
    .d1(q_32_25),
    .q(q_33_25)
  );
  

  flop_with_mux u_33_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_25),
    .d1(q_32_26),
    .q(q_33_26)
  );
  

  flop_with_mux u_33_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_26),
    .d1(q_32_27),
    .q(q_33_27)
  );
  

  flop_with_mux u_33_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_27),
    .d1(q_32_28),
    .q(q_33_28)
  );
  

  flop_with_mux u_33_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_28),
    .d1(q_32_29),
    .q(q_33_29)
  );
  

  flop_with_mux u_33_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_29),
    .d1(q_32_30),
    .q(q_33_30)
  );
  

  flop_with_mux u_33_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_30),
    .d1(q_32_31),
    .q(q_33_31)
  );
  

  flop_with_mux u_33_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_31),
    .d1(q_32_32),
    .q(q_33_32)
  );
  

  flop_with_mux u_33_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_32),
    .d1(q_32_33),
    .q(q_33_33)
  );
  

  flop_with_mux u_33_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_33),
    .d1(q_32_34),
    .q(q_33_34)
  );
  

  flop_with_mux u_33_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_34),
    .d1(q_32_35),
    .q(q_33_35)
  );
  

  flop_with_mux u_33_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_35),
    .d1(q_32_36),
    .q(q_33_36)
  );
  

  flop_with_mux u_33_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_36),
    .d1(q_32_37),
    .q(q_33_37)
  );
  

  flop_with_mux u_33_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_37),
    .d1(q_32_38),
    .q(q_33_38)
  );
  

  flop_with_mux u_33_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_38),
    .d1(q_32_39),
    .q(q_33_39)
  );
  

  flop_with_mux u_34_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_minus1),
    .d1(q_33_0),
    .q(q_34_0)
  );
  

  flop_with_mux u_34_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_0),
    .d1(q_33_1),
    .q(q_34_1)
  );
  

  flop_with_mux u_34_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_1),
    .d1(q_33_2),
    .q(q_34_2)
  );
  

  flop_with_mux u_34_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_2),
    .d1(q_33_3),
    .q(q_34_3)
  );
  

  flop_with_mux u_34_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_3),
    .d1(q_33_4),
    .q(q_34_4)
  );
  

  flop_with_mux u_34_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_4),
    .d1(q_33_5),
    .q(q_34_5)
  );
  

  flop_with_mux u_34_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_5),
    .d1(q_33_6),
    .q(q_34_6)
  );
  

  flop_with_mux u_34_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_6),
    .d1(q_33_7),
    .q(q_34_7)
  );
  

  flop_with_mux u_34_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_7),
    .d1(q_33_8),
    .q(q_34_8)
  );
  

  flop_with_mux u_34_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_8),
    .d1(q_33_9),
    .q(q_34_9)
  );
  

  flop_with_mux u_34_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_9),
    .d1(q_33_10),
    .q(q_34_10)
  );
  

  flop_with_mux u_34_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_10),
    .d1(q_33_11),
    .q(q_34_11)
  );
  

  flop_with_mux u_34_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_11),
    .d1(q_33_12),
    .q(q_34_12)
  );
  

  flop_with_mux u_34_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_12),
    .d1(q_33_13),
    .q(q_34_13)
  );
  

  flop_with_mux u_34_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_13),
    .d1(q_33_14),
    .q(q_34_14)
  );
  

  flop_with_mux u_34_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_14),
    .d1(q_33_15),
    .q(q_34_15)
  );
  

  flop_with_mux u_34_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_15),
    .d1(q_33_16),
    .q(q_34_16)
  );
  

  flop_with_mux u_34_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_16),
    .d1(q_33_17),
    .q(q_34_17)
  );
  

  flop_with_mux u_34_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_17),
    .d1(q_33_18),
    .q(q_34_18)
  );
  

  flop_with_mux u_34_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_18),
    .d1(q_33_19),
    .q(q_34_19)
  );
  

  flop_with_mux u_34_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_19),
    .d1(q_33_20),
    .q(q_34_20)
  );
  

  flop_with_mux u_34_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_20),
    .d1(q_33_21),
    .q(q_34_21)
  );
  

  flop_with_mux u_34_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_21),
    .d1(q_33_22),
    .q(q_34_22)
  );
  

  flop_with_mux u_34_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_22),
    .d1(q_33_23),
    .q(q_34_23)
  );
  

  flop_with_mux u_34_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_23),
    .d1(q_33_24),
    .q(q_34_24)
  );
  

  flop_with_mux u_34_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_24),
    .d1(q_33_25),
    .q(q_34_25)
  );
  

  flop_with_mux u_34_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_25),
    .d1(q_33_26),
    .q(q_34_26)
  );
  

  flop_with_mux u_34_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_26),
    .d1(q_33_27),
    .q(q_34_27)
  );
  

  flop_with_mux u_34_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_27),
    .d1(q_33_28),
    .q(q_34_28)
  );
  

  flop_with_mux u_34_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_28),
    .d1(q_33_29),
    .q(q_34_29)
  );
  

  flop_with_mux u_34_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_29),
    .d1(q_33_30),
    .q(q_34_30)
  );
  

  flop_with_mux u_34_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_30),
    .d1(q_33_31),
    .q(q_34_31)
  );
  

  flop_with_mux u_34_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_31),
    .d1(q_33_32),
    .q(q_34_32)
  );
  

  flop_with_mux u_34_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_32),
    .d1(q_33_33),
    .q(q_34_33)
  );
  

  flop_with_mux u_34_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_33),
    .d1(q_33_34),
    .q(q_34_34)
  );
  

  flop_with_mux u_34_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_34),
    .d1(q_33_35),
    .q(q_34_35)
  );
  

  flop_with_mux u_34_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_35),
    .d1(q_33_36),
    .q(q_34_36)
  );
  

  flop_with_mux u_34_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_36),
    .d1(q_33_37),
    .q(q_34_37)
  );
  

  flop_with_mux u_34_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_37),
    .d1(q_33_38),
    .q(q_34_38)
  );
  

  flop_with_mux u_34_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_38),
    .d1(q_33_39),
    .q(q_34_39)
  );
  

  flop_with_mux u_35_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_minus1),
    .d1(q_34_0),
    .q(q_35_0)
  );
  

  flop_with_mux u_35_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_0),
    .d1(q_34_1),
    .q(q_35_1)
  );
  

  flop_with_mux u_35_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_1),
    .d1(q_34_2),
    .q(q_35_2)
  );
  

  flop_with_mux u_35_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_2),
    .d1(q_34_3),
    .q(q_35_3)
  );
  

  flop_with_mux u_35_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_3),
    .d1(q_34_4),
    .q(q_35_4)
  );
  

  flop_with_mux u_35_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_4),
    .d1(q_34_5),
    .q(q_35_5)
  );
  

  flop_with_mux u_35_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_5),
    .d1(q_34_6),
    .q(q_35_6)
  );
  

  flop_with_mux u_35_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_6),
    .d1(q_34_7),
    .q(q_35_7)
  );
  

  flop_with_mux u_35_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_7),
    .d1(q_34_8),
    .q(q_35_8)
  );
  

  flop_with_mux u_35_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_8),
    .d1(q_34_9),
    .q(q_35_9)
  );
  

  flop_with_mux u_35_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_9),
    .d1(q_34_10),
    .q(q_35_10)
  );
  

  flop_with_mux u_35_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_10),
    .d1(q_34_11),
    .q(q_35_11)
  );
  

  flop_with_mux u_35_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_11),
    .d1(q_34_12),
    .q(q_35_12)
  );
  

  flop_with_mux u_35_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_12),
    .d1(q_34_13),
    .q(q_35_13)
  );
  

  flop_with_mux u_35_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_13),
    .d1(q_34_14),
    .q(q_35_14)
  );
  

  flop_with_mux u_35_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_14),
    .d1(q_34_15),
    .q(q_35_15)
  );
  

  flop_with_mux u_35_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_15),
    .d1(q_34_16),
    .q(q_35_16)
  );
  

  flop_with_mux u_35_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_16),
    .d1(q_34_17),
    .q(q_35_17)
  );
  

  flop_with_mux u_35_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_17),
    .d1(q_34_18),
    .q(q_35_18)
  );
  

  flop_with_mux u_35_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_18),
    .d1(q_34_19),
    .q(q_35_19)
  );
  

  flop_with_mux u_35_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_19),
    .d1(q_34_20),
    .q(q_35_20)
  );
  

  flop_with_mux u_35_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_20),
    .d1(q_34_21),
    .q(q_35_21)
  );
  

  flop_with_mux u_35_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_21),
    .d1(q_34_22),
    .q(q_35_22)
  );
  

  flop_with_mux u_35_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_22),
    .d1(q_34_23),
    .q(q_35_23)
  );
  

  flop_with_mux u_35_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_23),
    .d1(q_34_24),
    .q(q_35_24)
  );
  

  flop_with_mux u_35_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_24),
    .d1(q_34_25),
    .q(q_35_25)
  );
  

  flop_with_mux u_35_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_25),
    .d1(q_34_26),
    .q(q_35_26)
  );
  

  flop_with_mux u_35_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_26),
    .d1(q_34_27),
    .q(q_35_27)
  );
  

  flop_with_mux u_35_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_27),
    .d1(q_34_28),
    .q(q_35_28)
  );
  

  flop_with_mux u_35_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_28),
    .d1(q_34_29),
    .q(q_35_29)
  );
  

  flop_with_mux u_35_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_29),
    .d1(q_34_30),
    .q(q_35_30)
  );
  

  flop_with_mux u_35_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_30),
    .d1(q_34_31),
    .q(q_35_31)
  );
  

  flop_with_mux u_35_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_31),
    .d1(q_34_32),
    .q(q_35_32)
  );
  

  flop_with_mux u_35_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_32),
    .d1(q_34_33),
    .q(q_35_33)
  );
  

  flop_with_mux u_35_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_33),
    .d1(q_34_34),
    .q(q_35_34)
  );
  

  flop_with_mux u_35_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_34),
    .d1(q_34_35),
    .q(q_35_35)
  );
  

  flop_with_mux u_35_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_35),
    .d1(q_34_36),
    .q(q_35_36)
  );
  

  flop_with_mux u_35_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_36),
    .d1(q_34_37),
    .q(q_35_37)
  );
  

  flop_with_mux u_35_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_37),
    .d1(q_34_38),
    .q(q_35_38)
  );
  

  flop_with_mux u_35_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_38),
    .d1(q_34_39),
    .q(q_35_39)
  );
  

  flop_with_mux u_36_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_minus1),
    .d1(q_35_0),
    .q(q_36_0)
  );
  

  flop_with_mux u_36_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_0),
    .d1(q_35_1),
    .q(q_36_1)
  );
  

  flop_with_mux u_36_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_1),
    .d1(q_35_2),
    .q(q_36_2)
  );
  

  flop_with_mux u_36_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_2),
    .d1(q_35_3),
    .q(q_36_3)
  );
  

  flop_with_mux u_36_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_3),
    .d1(q_35_4),
    .q(q_36_4)
  );
  

  flop_with_mux u_36_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_4),
    .d1(q_35_5),
    .q(q_36_5)
  );
  

  flop_with_mux u_36_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_5),
    .d1(q_35_6),
    .q(q_36_6)
  );
  

  flop_with_mux u_36_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_6),
    .d1(q_35_7),
    .q(q_36_7)
  );
  

  flop_with_mux u_36_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_7),
    .d1(q_35_8),
    .q(q_36_8)
  );
  

  flop_with_mux u_36_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_8),
    .d1(q_35_9),
    .q(q_36_9)
  );
  

  flop_with_mux u_36_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_9),
    .d1(q_35_10),
    .q(q_36_10)
  );
  

  flop_with_mux u_36_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_10),
    .d1(q_35_11),
    .q(q_36_11)
  );
  

  flop_with_mux u_36_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_11),
    .d1(q_35_12),
    .q(q_36_12)
  );
  

  flop_with_mux u_36_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_12),
    .d1(q_35_13),
    .q(q_36_13)
  );
  

  flop_with_mux u_36_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_13),
    .d1(q_35_14),
    .q(q_36_14)
  );
  

  flop_with_mux u_36_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_14),
    .d1(q_35_15),
    .q(q_36_15)
  );
  

  flop_with_mux u_36_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_15),
    .d1(q_35_16),
    .q(q_36_16)
  );
  

  flop_with_mux u_36_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_16),
    .d1(q_35_17),
    .q(q_36_17)
  );
  

  flop_with_mux u_36_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_17),
    .d1(q_35_18),
    .q(q_36_18)
  );
  

  flop_with_mux u_36_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_18),
    .d1(q_35_19),
    .q(q_36_19)
  );
  

  flop_with_mux u_36_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_19),
    .d1(q_35_20),
    .q(q_36_20)
  );
  

  flop_with_mux u_36_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_20),
    .d1(q_35_21),
    .q(q_36_21)
  );
  

  flop_with_mux u_36_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_21),
    .d1(q_35_22),
    .q(q_36_22)
  );
  

  flop_with_mux u_36_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_22),
    .d1(q_35_23),
    .q(q_36_23)
  );
  

  flop_with_mux u_36_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_23),
    .d1(q_35_24),
    .q(q_36_24)
  );
  

  flop_with_mux u_36_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_24),
    .d1(q_35_25),
    .q(q_36_25)
  );
  

  flop_with_mux u_36_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_25),
    .d1(q_35_26),
    .q(q_36_26)
  );
  

  flop_with_mux u_36_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_26),
    .d1(q_35_27),
    .q(q_36_27)
  );
  

  flop_with_mux u_36_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_27),
    .d1(q_35_28),
    .q(q_36_28)
  );
  

  flop_with_mux u_36_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_28),
    .d1(q_35_29),
    .q(q_36_29)
  );
  

  flop_with_mux u_36_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_29),
    .d1(q_35_30),
    .q(q_36_30)
  );
  

  flop_with_mux u_36_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_30),
    .d1(q_35_31),
    .q(q_36_31)
  );
  

  flop_with_mux u_36_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_31),
    .d1(q_35_32),
    .q(q_36_32)
  );
  

  flop_with_mux u_36_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_32),
    .d1(q_35_33),
    .q(q_36_33)
  );
  

  flop_with_mux u_36_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_33),
    .d1(q_35_34),
    .q(q_36_34)
  );
  

  flop_with_mux u_36_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_34),
    .d1(q_35_35),
    .q(q_36_35)
  );
  

  flop_with_mux u_36_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_35),
    .d1(q_35_36),
    .q(q_36_36)
  );
  

  flop_with_mux u_36_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_36),
    .d1(q_35_37),
    .q(q_36_37)
  );
  

  flop_with_mux u_36_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_37),
    .d1(q_35_38),
    .q(q_36_38)
  );
  

  flop_with_mux u_36_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_38),
    .d1(q_35_39),
    .q(q_36_39)
  );
  

  flop_with_mux u_37_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_minus1),
    .d1(q_36_0),
    .q(q_37_0)
  );
  

  flop_with_mux u_37_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_0),
    .d1(q_36_1),
    .q(q_37_1)
  );
  

  flop_with_mux u_37_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_1),
    .d1(q_36_2),
    .q(q_37_2)
  );
  

  flop_with_mux u_37_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_2),
    .d1(q_36_3),
    .q(q_37_3)
  );
  

  flop_with_mux u_37_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_3),
    .d1(q_36_4),
    .q(q_37_4)
  );
  

  flop_with_mux u_37_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_4),
    .d1(q_36_5),
    .q(q_37_5)
  );
  

  flop_with_mux u_37_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_5),
    .d1(q_36_6),
    .q(q_37_6)
  );
  

  flop_with_mux u_37_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_6),
    .d1(q_36_7),
    .q(q_37_7)
  );
  

  flop_with_mux u_37_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_7),
    .d1(q_36_8),
    .q(q_37_8)
  );
  

  flop_with_mux u_37_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_8),
    .d1(q_36_9),
    .q(q_37_9)
  );
  

  flop_with_mux u_37_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_9),
    .d1(q_36_10),
    .q(q_37_10)
  );
  

  flop_with_mux u_37_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_10),
    .d1(q_36_11),
    .q(q_37_11)
  );
  

  flop_with_mux u_37_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_11),
    .d1(q_36_12),
    .q(q_37_12)
  );
  

  flop_with_mux u_37_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_12),
    .d1(q_36_13),
    .q(q_37_13)
  );
  

  flop_with_mux u_37_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_13),
    .d1(q_36_14),
    .q(q_37_14)
  );
  

  flop_with_mux u_37_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_14),
    .d1(q_36_15),
    .q(q_37_15)
  );
  

  flop_with_mux u_37_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_15),
    .d1(q_36_16),
    .q(q_37_16)
  );
  

  flop_with_mux u_37_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_16),
    .d1(q_36_17),
    .q(q_37_17)
  );
  

  flop_with_mux u_37_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_17),
    .d1(q_36_18),
    .q(q_37_18)
  );
  

  flop_with_mux u_37_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_18),
    .d1(q_36_19),
    .q(q_37_19)
  );
  

  flop_with_mux u_37_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_19),
    .d1(q_36_20),
    .q(q_37_20)
  );
  

  flop_with_mux u_37_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_20),
    .d1(q_36_21),
    .q(q_37_21)
  );
  

  flop_with_mux u_37_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_21),
    .d1(q_36_22),
    .q(q_37_22)
  );
  

  flop_with_mux u_37_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_22),
    .d1(q_36_23),
    .q(q_37_23)
  );
  

  flop_with_mux u_37_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_23),
    .d1(q_36_24),
    .q(q_37_24)
  );
  

  flop_with_mux u_37_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_24),
    .d1(q_36_25),
    .q(q_37_25)
  );
  

  flop_with_mux u_37_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_25),
    .d1(q_36_26),
    .q(q_37_26)
  );
  

  flop_with_mux u_37_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_26),
    .d1(q_36_27),
    .q(q_37_27)
  );
  

  flop_with_mux u_37_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_27),
    .d1(q_36_28),
    .q(q_37_28)
  );
  

  flop_with_mux u_37_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_28),
    .d1(q_36_29),
    .q(q_37_29)
  );
  

  flop_with_mux u_37_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_29),
    .d1(q_36_30),
    .q(q_37_30)
  );
  

  flop_with_mux u_37_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_30),
    .d1(q_36_31),
    .q(q_37_31)
  );
  

  flop_with_mux u_37_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_31),
    .d1(q_36_32),
    .q(q_37_32)
  );
  

  flop_with_mux u_37_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_32),
    .d1(q_36_33),
    .q(q_37_33)
  );
  

  flop_with_mux u_37_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_33),
    .d1(q_36_34),
    .q(q_37_34)
  );
  

  flop_with_mux u_37_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_34),
    .d1(q_36_35),
    .q(q_37_35)
  );
  

  flop_with_mux u_37_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_35),
    .d1(q_36_36),
    .q(q_37_36)
  );
  

  flop_with_mux u_37_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_36),
    .d1(q_36_37),
    .q(q_37_37)
  );
  

  flop_with_mux u_37_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_37),
    .d1(q_36_38),
    .q(q_37_38)
  );
  

  flop_with_mux u_37_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_38),
    .d1(q_36_39),
    .q(q_37_39)
  );
  

  flop_with_mux u_38_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_minus1),
    .d1(q_37_0),
    .q(q_38_0)
  );
  

  flop_with_mux u_38_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_0),
    .d1(q_37_1),
    .q(q_38_1)
  );
  

  flop_with_mux u_38_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_1),
    .d1(q_37_2),
    .q(q_38_2)
  );
  

  flop_with_mux u_38_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_2),
    .d1(q_37_3),
    .q(q_38_3)
  );
  

  flop_with_mux u_38_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_3),
    .d1(q_37_4),
    .q(q_38_4)
  );
  

  flop_with_mux u_38_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_4),
    .d1(q_37_5),
    .q(q_38_5)
  );
  

  flop_with_mux u_38_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_5),
    .d1(q_37_6),
    .q(q_38_6)
  );
  

  flop_with_mux u_38_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_6),
    .d1(q_37_7),
    .q(q_38_7)
  );
  

  flop_with_mux u_38_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_7),
    .d1(q_37_8),
    .q(q_38_8)
  );
  

  flop_with_mux u_38_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_8),
    .d1(q_37_9),
    .q(q_38_9)
  );
  

  flop_with_mux u_38_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_9),
    .d1(q_37_10),
    .q(q_38_10)
  );
  

  flop_with_mux u_38_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_10),
    .d1(q_37_11),
    .q(q_38_11)
  );
  

  flop_with_mux u_38_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_11),
    .d1(q_37_12),
    .q(q_38_12)
  );
  

  flop_with_mux u_38_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_12),
    .d1(q_37_13),
    .q(q_38_13)
  );
  

  flop_with_mux u_38_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_13),
    .d1(q_37_14),
    .q(q_38_14)
  );
  

  flop_with_mux u_38_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_14),
    .d1(q_37_15),
    .q(q_38_15)
  );
  

  flop_with_mux u_38_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_15),
    .d1(q_37_16),
    .q(q_38_16)
  );
  

  flop_with_mux u_38_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_16),
    .d1(q_37_17),
    .q(q_38_17)
  );
  

  flop_with_mux u_38_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_17),
    .d1(q_37_18),
    .q(q_38_18)
  );
  

  flop_with_mux u_38_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_18),
    .d1(q_37_19),
    .q(q_38_19)
  );
  

  flop_with_mux u_38_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_19),
    .d1(q_37_20),
    .q(q_38_20)
  );
  

  flop_with_mux u_38_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_20),
    .d1(q_37_21),
    .q(q_38_21)
  );
  

  flop_with_mux u_38_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_21),
    .d1(q_37_22),
    .q(q_38_22)
  );
  

  flop_with_mux u_38_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_22),
    .d1(q_37_23),
    .q(q_38_23)
  );
  

  flop_with_mux u_38_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_23),
    .d1(q_37_24),
    .q(q_38_24)
  );
  

  flop_with_mux u_38_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_24),
    .d1(q_37_25),
    .q(q_38_25)
  );
  

  flop_with_mux u_38_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_25),
    .d1(q_37_26),
    .q(q_38_26)
  );
  

  flop_with_mux u_38_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_26),
    .d1(q_37_27),
    .q(q_38_27)
  );
  

  flop_with_mux u_38_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_27),
    .d1(q_37_28),
    .q(q_38_28)
  );
  

  flop_with_mux u_38_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_28),
    .d1(q_37_29),
    .q(q_38_29)
  );
  

  flop_with_mux u_38_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_29),
    .d1(q_37_30),
    .q(q_38_30)
  );
  

  flop_with_mux u_38_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_30),
    .d1(q_37_31),
    .q(q_38_31)
  );
  

  flop_with_mux u_38_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_31),
    .d1(q_37_32),
    .q(q_38_32)
  );
  

  flop_with_mux u_38_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_32),
    .d1(q_37_33),
    .q(q_38_33)
  );
  

  flop_with_mux u_38_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_33),
    .d1(q_37_34),
    .q(q_38_34)
  );
  

  flop_with_mux u_38_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_34),
    .d1(q_37_35),
    .q(q_38_35)
  );
  

  flop_with_mux u_38_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_35),
    .d1(q_37_36),
    .q(q_38_36)
  );
  

  flop_with_mux u_38_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_36),
    .d1(q_37_37),
    .q(q_38_37)
  );
  

  flop_with_mux u_38_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_37),
    .d1(q_37_38),
    .q(q_38_38)
  );
  

  flop_with_mux u_38_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_38),
    .d1(q_37_39),
    .q(q_38_39)
  );
  

  flop_with_mux u_39_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_minus1),
    .d1(q_38_0),
    .q(q_39_0)
  );
  

  flop_with_mux u_39_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_0),
    .d1(q_38_1),
    .q(q_39_1)
  );
  

  flop_with_mux u_39_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_1),
    .d1(q_38_2),
    .q(q_39_2)
  );
  

  flop_with_mux u_39_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_2),
    .d1(q_38_3),
    .q(q_39_3)
  );
  

  flop_with_mux u_39_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_3),
    .d1(q_38_4),
    .q(q_39_4)
  );
  

  flop_with_mux u_39_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_4),
    .d1(q_38_5),
    .q(q_39_5)
  );
  

  flop_with_mux u_39_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_5),
    .d1(q_38_6),
    .q(q_39_6)
  );
  

  flop_with_mux u_39_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_6),
    .d1(q_38_7),
    .q(q_39_7)
  );
  

  flop_with_mux u_39_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_7),
    .d1(q_38_8),
    .q(q_39_8)
  );
  

  flop_with_mux u_39_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_8),
    .d1(q_38_9),
    .q(q_39_9)
  );
  

  flop_with_mux u_39_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_9),
    .d1(q_38_10),
    .q(q_39_10)
  );
  

  flop_with_mux u_39_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_10),
    .d1(q_38_11),
    .q(q_39_11)
  );
  

  flop_with_mux u_39_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_11),
    .d1(q_38_12),
    .q(q_39_12)
  );
  

  flop_with_mux u_39_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_12),
    .d1(q_38_13),
    .q(q_39_13)
  );
  

  flop_with_mux u_39_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_13),
    .d1(q_38_14),
    .q(q_39_14)
  );
  

  flop_with_mux u_39_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_14),
    .d1(q_38_15),
    .q(q_39_15)
  );
  

  flop_with_mux u_39_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_15),
    .d1(q_38_16),
    .q(q_39_16)
  );
  

  flop_with_mux u_39_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_16),
    .d1(q_38_17),
    .q(q_39_17)
  );
  

  flop_with_mux u_39_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_17),
    .d1(q_38_18),
    .q(q_39_18)
  );
  

  flop_with_mux u_39_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_18),
    .d1(q_38_19),
    .q(q_39_19)
  );
  

  flop_with_mux u_39_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_19),
    .d1(q_38_20),
    .q(q_39_20)
  );
  

  flop_with_mux u_39_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_20),
    .d1(q_38_21),
    .q(q_39_21)
  );
  

  flop_with_mux u_39_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_21),
    .d1(q_38_22),
    .q(q_39_22)
  );
  

  flop_with_mux u_39_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_22),
    .d1(q_38_23),
    .q(q_39_23)
  );
  

  flop_with_mux u_39_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_23),
    .d1(q_38_24),
    .q(q_39_24)
  );
  

  flop_with_mux u_39_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_24),
    .d1(q_38_25),
    .q(q_39_25)
  );
  

  flop_with_mux u_39_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_25),
    .d1(q_38_26),
    .q(q_39_26)
  );
  

  flop_with_mux u_39_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_26),
    .d1(q_38_27),
    .q(q_39_27)
  );
  

  flop_with_mux u_39_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_27),
    .d1(q_38_28),
    .q(q_39_28)
  );
  

  flop_with_mux u_39_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_28),
    .d1(q_38_29),
    .q(q_39_29)
  );
  

  flop_with_mux u_39_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_29),
    .d1(q_38_30),
    .q(q_39_30)
  );
  

  flop_with_mux u_39_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_30),
    .d1(q_38_31),
    .q(q_39_31)
  );
  

  flop_with_mux u_39_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_31),
    .d1(q_38_32),
    .q(q_39_32)
  );
  

  flop_with_mux u_39_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_32),
    .d1(q_38_33),
    .q(q_39_33)
  );
  

  flop_with_mux u_39_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_33),
    .d1(q_38_34),
    .q(q_39_34)
  );
  

  flop_with_mux u_39_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_34),
    .d1(q_38_35),
    .q(q_39_35)
  );
  

  flop_with_mux u_39_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_35),
    .d1(q_38_36),
    .q(q_39_36)
  );
  

  flop_with_mux u_39_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_36),
    .d1(q_38_37),
    .q(q_39_37)
  );
  

  flop_with_mux u_39_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_37),
    .d1(q_38_38),
    .q(q_39_38)
  );
  

  flop_with_mux u_39_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_38),
    .d1(q_38_39),
    .q(q_39_39)
  );
  
endmodule

  module pong_buffer (
  input [40-1:0] data_in,
  output [40-1:0] data_out,
  input load_unload, //0 for load (left to right), 1 for unload (top to bottom)
  input valid,
  input clk);

  wire [40-1:0] data_out_internal;
  assign data_out = data_out_internal & {40{load_unload}};
  
wire q_0_0;
wire q_0_1;
wire q_0_2;
wire q_0_3;
wire q_0_4;
wire q_0_5;
wire q_0_6;
wire q_0_7;
wire q_0_8;
wire q_0_9;
wire q_0_10;
wire q_0_11;
wire q_0_12;
wire q_0_13;
wire q_0_14;
wire q_0_15;
wire q_0_16;
wire q_0_17;
wire q_0_18;
wire q_0_19;
wire q_0_20;
wire q_0_21;
wire q_0_22;
wire q_0_23;
wire q_0_24;
wire q_0_25;
wire q_0_26;
wire q_0_27;
wire q_0_28;
wire q_0_29;
wire q_0_30;
wire q_0_31;
wire q_0_32;
wire q_0_33;
wire q_0_34;
wire q_0_35;
wire q_0_36;
wire q_0_37;
wire q_0_38;
wire q_0_39;
wire q_1_0;
wire q_1_1;
wire q_1_2;
wire q_1_3;
wire q_1_4;
wire q_1_5;
wire q_1_6;
wire q_1_7;
wire q_1_8;
wire q_1_9;
wire q_1_10;
wire q_1_11;
wire q_1_12;
wire q_1_13;
wire q_1_14;
wire q_1_15;
wire q_1_16;
wire q_1_17;
wire q_1_18;
wire q_1_19;
wire q_1_20;
wire q_1_21;
wire q_1_22;
wire q_1_23;
wire q_1_24;
wire q_1_25;
wire q_1_26;
wire q_1_27;
wire q_1_28;
wire q_1_29;
wire q_1_30;
wire q_1_31;
wire q_1_32;
wire q_1_33;
wire q_1_34;
wire q_1_35;
wire q_1_36;
wire q_1_37;
wire q_1_38;
wire q_1_39;
wire q_2_0;
wire q_2_1;
wire q_2_2;
wire q_2_3;
wire q_2_4;
wire q_2_5;
wire q_2_6;
wire q_2_7;
wire q_2_8;
wire q_2_9;
wire q_2_10;
wire q_2_11;
wire q_2_12;
wire q_2_13;
wire q_2_14;
wire q_2_15;
wire q_2_16;
wire q_2_17;
wire q_2_18;
wire q_2_19;
wire q_2_20;
wire q_2_21;
wire q_2_22;
wire q_2_23;
wire q_2_24;
wire q_2_25;
wire q_2_26;
wire q_2_27;
wire q_2_28;
wire q_2_29;
wire q_2_30;
wire q_2_31;
wire q_2_32;
wire q_2_33;
wire q_2_34;
wire q_2_35;
wire q_2_36;
wire q_2_37;
wire q_2_38;
wire q_2_39;
wire q_3_0;
wire q_3_1;
wire q_3_2;
wire q_3_3;
wire q_3_4;
wire q_3_5;
wire q_3_6;
wire q_3_7;
wire q_3_8;
wire q_3_9;
wire q_3_10;
wire q_3_11;
wire q_3_12;
wire q_3_13;
wire q_3_14;
wire q_3_15;
wire q_3_16;
wire q_3_17;
wire q_3_18;
wire q_3_19;
wire q_3_20;
wire q_3_21;
wire q_3_22;
wire q_3_23;
wire q_3_24;
wire q_3_25;
wire q_3_26;
wire q_3_27;
wire q_3_28;
wire q_3_29;
wire q_3_30;
wire q_3_31;
wire q_3_32;
wire q_3_33;
wire q_3_34;
wire q_3_35;
wire q_3_36;
wire q_3_37;
wire q_3_38;
wire q_3_39;
wire q_4_0;
wire q_4_1;
wire q_4_2;
wire q_4_3;
wire q_4_4;
wire q_4_5;
wire q_4_6;
wire q_4_7;
wire q_4_8;
wire q_4_9;
wire q_4_10;
wire q_4_11;
wire q_4_12;
wire q_4_13;
wire q_4_14;
wire q_4_15;
wire q_4_16;
wire q_4_17;
wire q_4_18;
wire q_4_19;
wire q_4_20;
wire q_4_21;
wire q_4_22;
wire q_4_23;
wire q_4_24;
wire q_4_25;
wire q_4_26;
wire q_4_27;
wire q_4_28;
wire q_4_29;
wire q_4_30;
wire q_4_31;
wire q_4_32;
wire q_4_33;
wire q_4_34;
wire q_4_35;
wire q_4_36;
wire q_4_37;
wire q_4_38;
wire q_4_39;
wire q_5_0;
wire q_5_1;
wire q_5_2;
wire q_5_3;
wire q_5_4;
wire q_5_5;
wire q_5_6;
wire q_5_7;
wire q_5_8;
wire q_5_9;
wire q_5_10;
wire q_5_11;
wire q_5_12;
wire q_5_13;
wire q_5_14;
wire q_5_15;
wire q_5_16;
wire q_5_17;
wire q_5_18;
wire q_5_19;
wire q_5_20;
wire q_5_21;
wire q_5_22;
wire q_5_23;
wire q_5_24;
wire q_5_25;
wire q_5_26;
wire q_5_27;
wire q_5_28;
wire q_5_29;
wire q_5_30;
wire q_5_31;
wire q_5_32;
wire q_5_33;
wire q_5_34;
wire q_5_35;
wire q_5_36;
wire q_5_37;
wire q_5_38;
wire q_5_39;
wire q_6_0;
wire q_6_1;
wire q_6_2;
wire q_6_3;
wire q_6_4;
wire q_6_5;
wire q_6_6;
wire q_6_7;
wire q_6_8;
wire q_6_9;
wire q_6_10;
wire q_6_11;
wire q_6_12;
wire q_6_13;
wire q_6_14;
wire q_6_15;
wire q_6_16;
wire q_6_17;
wire q_6_18;
wire q_6_19;
wire q_6_20;
wire q_6_21;
wire q_6_22;
wire q_6_23;
wire q_6_24;
wire q_6_25;
wire q_6_26;
wire q_6_27;
wire q_6_28;
wire q_6_29;
wire q_6_30;
wire q_6_31;
wire q_6_32;
wire q_6_33;
wire q_6_34;
wire q_6_35;
wire q_6_36;
wire q_6_37;
wire q_6_38;
wire q_6_39;
wire q_7_0;
wire q_7_1;
wire q_7_2;
wire q_7_3;
wire q_7_4;
wire q_7_5;
wire q_7_6;
wire q_7_7;
wire q_7_8;
wire q_7_9;
wire q_7_10;
wire q_7_11;
wire q_7_12;
wire q_7_13;
wire q_7_14;
wire q_7_15;
wire q_7_16;
wire q_7_17;
wire q_7_18;
wire q_7_19;
wire q_7_20;
wire q_7_21;
wire q_7_22;
wire q_7_23;
wire q_7_24;
wire q_7_25;
wire q_7_26;
wire q_7_27;
wire q_7_28;
wire q_7_29;
wire q_7_30;
wire q_7_31;
wire q_7_32;
wire q_7_33;
wire q_7_34;
wire q_7_35;
wire q_7_36;
wire q_7_37;
wire q_7_38;
wire q_7_39;
wire q_8_0;
wire q_8_1;
wire q_8_2;
wire q_8_3;
wire q_8_4;
wire q_8_5;
wire q_8_6;
wire q_8_7;
wire q_8_8;
wire q_8_9;
wire q_8_10;
wire q_8_11;
wire q_8_12;
wire q_8_13;
wire q_8_14;
wire q_8_15;
wire q_8_16;
wire q_8_17;
wire q_8_18;
wire q_8_19;
wire q_8_20;
wire q_8_21;
wire q_8_22;
wire q_8_23;
wire q_8_24;
wire q_8_25;
wire q_8_26;
wire q_8_27;
wire q_8_28;
wire q_8_29;
wire q_8_30;
wire q_8_31;
wire q_8_32;
wire q_8_33;
wire q_8_34;
wire q_8_35;
wire q_8_36;
wire q_8_37;
wire q_8_38;
wire q_8_39;
wire q_9_0;
wire q_9_1;
wire q_9_2;
wire q_9_3;
wire q_9_4;
wire q_9_5;
wire q_9_6;
wire q_9_7;
wire q_9_8;
wire q_9_9;
wire q_9_10;
wire q_9_11;
wire q_9_12;
wire q_9_13;
wire q_9_14;
wire q_9_15;
wire q_9_16;
wire q_9_17;
wire q_9_18;
wire q_9_19;
wire q_9_20;
wire q_9_21;
wire q_9_22;
wire q_9_23;
wire q_9_24;
wire q_9_25;
wire q_9_26;
wire q_9_27;
wire q_9_28;
wire q_9_29;
wire q_9_30;
wire q_9_31;
wire q_9_32;
wire q_9_33;
wire q_9_34;
wire q_9_35;
wire q_9_36;
wire q_9_37;
wire q_9_38;
wire q_9_39;
wire q_10_0;
wire q_10_1;
wire q_10_2;
wire q_10_3;
wire q_10_4;
wire q_10_5;
wire q_10_6;
wire q_10_7;
wire q_10_8;
wire q_10_9;
wire q_10_10;
wire q_10_11;
wire q_10_12;
wire q_10_13;
wire q_10_14;
wire q_10_15;
wire q_10_16;
wire q_10_17;
wire q_10_18;
wire q_10_19;
wire q_10_20;
wire q_10_21;
wire q_10_22;
wire q_10_23;
wire q_10_24;
wire q_10_25;
wire q_10_26;
wire q_10_27;
wire q_10_28;
wire q_10_29;
wire q_10_30;
wire q_10_31;
wire q_10_32;
wire q_10_33;
wire q_10_34;
wire q_10_35;
wire q_10_36;
wire q_10_37;
wire q_10_38;
wire q_10_39;
wire q_11_0;
wire q_11_1;
wire q_11_2;
wire q_11_3;
wire q_11_4;
wire q_11_5;
wire q_11_6;
wire q_11_7;
wire q_11_8;
wire q_11_9;
wire q_11_10;
wire q_11_11;
wire q_11_12;
wire q_11_13;
wire q_11_14;
wire q_11_15;
wire q_11_16;
wire q_11_17;
wire q_11_18;
wire q_11_19;
wire q_11_20;
wire q_11_21;
wire q_11_22;
wire q_11_23;
wire q_11_24;
wire q_11_25;
wire q_11_26;
wire q_11_27;
wire q_11_28;
wire q_11_29;
wire q_11_30;
wire q_11_31;
wire q_11_32;
wire q_11_33;
wire q_11_34;
wire q_11_35;
wire q_11_36;
wire q_11_37;
wire q_11_38;
wire q_11_39;
wire q_12_0;
wire q_12_1;
wire q_12_2;
wire q_12_3;
wire q_12_4;
wire q_12_5;
wire q_12_6;
wire q_12_7;
wire q_12_8;
wire q_12_9;
wire q_12_10;
wire q_12_11;
wire q_12_12;
wire q_12_13;
wire q_12_14;
wire q_12_15;
wire q_12_16;
wire q_12_17;
wire q_12_18;
wire q_12_19;
wire q_12_20;
wire q_12_21;
wire q_12_22;
wire q_12_23;
wire q_12_24;
wire q_12_25;
wire q_12_26;
wire q_12_27;
wire q_12_28;
wire q_12_29;
wire q_12_30;
wire q_12_31;
wire q_12_32;
wire q_12_33;
wire q_12_34;
wire q_12_35;
wire q_12_36;
wire q_12_37;
wire q_12_38;
wire q_12_39;
wire q_13_0;
wire q_13_1;
wire q_13_2;
wire q_13_3;
wire q_13_4;
wire q_13_5;
wire q_13_6;
wire q_13_7;
wire q_13_8;
wire q_13_9;
wire q_13_10;
wire q_13_11;
wire q_13_12;
wire q_13_13;
wire q_13_14;
wire q_13_15;
wire q_13_16;
wire q_13_17;
wire q_13_18;
wire q_13_19;
wire q_13_20;
wire q_13_21;
wire q_13_22;
wire q_13_23;
wire q_13_24;
wire q_13_25;
wire q_13_26;
wire q_13_27;
wire q_13_28;
wire q_13_29;
wire q_13_30;
wire q_13_31;
wire q_13_32;
wire q_13_33;
wire q_13_34;
wire q_13_35;
wire q_13_36;
wire q_13_37;
wire q_13_38;
wire q_13_39;
wire q_14_0;
wire q_14_1;
wire q_14_2;
wire q_14_3;
wire q_14_4;
wire q_14_5;
wire q_14_6;
wire q_14_7;
wire q_14_8;
wire q_14_9;
wire q_14_10;
wire q_14_11;
wire q_14_12;
wire q_14_13;
wire q_14_14;
wire q_14_15;
wire q_14_16;
wire q_14_17;
wire q_14_18;
wire q_14_19;
wire q_14_20;
wire q_14_21;
wire q_14_22;
wire q_14_23;
wire q_14_24;
wire q_14_25;
wire q_14_26;
wire q_14_27;
wire q_14_28;
wire q_14_29;
wire q_14_30;
wire q_14_31;
wire q_14_32;
wire q_14_33;
wire q_14_34;
wire q_14_35;
wire q_14_36;
wire q_14_37;
wire q_14_38;
wire q_14_39;
wire q_15_0;
wire q_15_1;
wire q_15_2;
wire q_15_3;
wire q_15_4;
wire q_15_5;
wire q_15_6;
wire q_15_7;
wire q_15_8;
wire q_15_9;
wire q_15_10;
wire q_15_11;
wire q_15_12;
wire q_15_13;
wire q_15_14;
wire q_15_15;
wire q_15_16;
wire q_15_17;
wire q_15_18;
wire q_15_19;
wire q_15_20;
wire q_15_21;
wire q_15_22;
wire q_15_23;
wire q_15_24;
wire q_15_25;
wire q_15_26;
wire q_15_27;
wire q_15_28;
wire q_15_29;
wire q_15_30;
wire q_15_31;
wire q_15_32;
wire q_15_33;
wire q_15_34;
wire q_15_35;
wire q_15_36;
wire q_15_37;
wire q_15_38;
wire q_15_39;
wire q_16_0;
wire q_16_1;
wire q_16_2;
wire q_16_3;
wire q_16_4;
wire q_16_5;
wire q_16_6;
wire q_16_7;
wire q_16_8;
wire q_16_9;
wire q_16_10;
wire q_16_11;
wire q_16_12;
wire q_16_13;
wire q_16_14;
wire q_16_15;
wire q_16_16;
wire q_16_17;
wire q_16_18;
wire q_16_19;
wire q_16_20;
wire q_16_21;
wire q_16_22;
wire q_16_23;
wire q_16_24;
wire q_16_25;
wire q_16_26;
wire q_16_27;
wire q_16_28;
wire q_16_29;
wire q_16_30;
wire q_16_31;
wire q_16_32;
wire q_16_33;
wire q_16_34;
wire q_16_35;
wire q_16_36;
wire q_16_37;
wire q_16_38;
wire q_16_39;
wire q_17_0;
wire q_17_1;
wire q_17_2;
wire q_17_3;
wire q_17_4;
wire q_17_5;
wire q_17_6;
wire q_17_7;
wire q_17_8;
wire q_17_9;
wire q_17_10;
wire q_17_11;
wire q_17_12;
wire q_17_13;
wire q_17_14;
wire q_17_15;
wire q_17_16;
wire q_17_17;
wire q_17_18;
wire q_17_19;
wire q_17_20;
wire q_17_21;
wire q_17_22;
wire q_17_23;
wire q_17_24;
wire q_17_25;
wire q_17_26;
wire q_17_27;
wire q_17_28;
wire q_17_29;
wire q_17_30;
wire q_17_31;
wire q_17_32;
wire q_17_33;
wire q_17_34;
wire q_17_35;
wire q_17_36;
wire q_17_37;
wire q_17_38;
wire q_17_39;
wire q_18_0;
wire q_18_1;
wire q_18_2;
wire q_18_3;
wire q_18_4;
wire q_18_5;
wire q_18_6;
wire q_18_7;
wire q_18_8;
wire q_18_9;
wire q_18_10;
wire q_18_11;
wire q_18_12;
wire q_18_13;
wire q_18_14;
wire q_18_15;
wire q_18_16;
wire q_18_17;
wire q_18_18;
wire q_18_19;
wire q_18_20;
wire q_18_21;
wire q_18_22;
wire q_18_23;
wire q_18_24;
wire q_18_25;
wire q_18_26;
wire q_18_27;
wire q_18_28;
wire q_18_29;
wire q_18_30;
wire q_18_31;
wire q_18_32;
wire q_18_33;
wire q_18_34;
wire q_18_35;
wire q_18_36;
wire q_18_37;
wire q_18_38;
wire q_18_39;
wire q_19_0;
wire q_19_1;
wire q_19_2;
wire q_19_3;
wire q_19_4;
wire q_19_5;
wire q_19_6;
wire q_19_7;
wire q_19_8;
wire q_19_9;
wire q_19_10;
wire q_19_11;
wire q_19_12;
wire q_19_13;
wire q_19_14;
wire q_19_15;
wire q_19_16;
wire q_19_17;
wire q_19_18;
wire q_19_19;
wire q_19_20;
wire q_19_21;
wire q_19_22;
wire q_19_23;
wire q_19_24;
wire q_19_25;
wire q_19_26;
wire q_19_27;
wire q_19_28;
wire q_19_29;
wire q_19_30;
wire q_19_31;
wire q_19_32;
wire q_19_33;
wire q_19_34;
wire q_19_35;
wire q_19_36;
wire q_19_37;
wire q_19_38;
wire q_19_39;
wire q_20_0;
wire q_20_1;
wire q_20_2;
wire q_20_3;
wire q_20_4;
wire q_20_5;
wire q_20_6;
wire q_20_7;
wire q_20_8;
wire q_20_9;
wire q_20_10;
wire q_20_11;
wire q_20_12;
wire q_20_13;
wire q_20_14;
wire q_20_15;
wire q_20_16;
wire q_20_17;
wire q_20_18;
wire q_20_19;
wire q_20_20;
wire q_20_21;
wire q_20_22;
wire q_20_23;
wire q_20_24;
wire q_20_25;
wire q_20_26;
wire q_20_27;
wire q_20_28;
wire q_20_29;
wire q_20_30;
wire q_20_31;
wire q_20_32;
wire q_20_33;
wire q_20_34;
wire q_20_35;
wire q_20_36;
wire q_20_37;
wire q_20_38;
wire q_20_39;
wire q_21_0;
wire q_21_1;
wire q_21_2;
wire q_21_3;
wire q_21_4;
wire q_21_5;
wire q_21_6;
wire q_21_7;
wire q_21_8;
wire q_21_9;
wire q_21_10;
wire q_21_11;
wire q_21_12;
wire q_21_13;
wire q_21_14;
wire q_21_15;
wire q_21_16;
wire q_21_17;
wire q_21_18;
wire q_21_19;
wire q_21_20;
wire q_21_21;
wire q_21_22;
wire q_21_23;
wire q_21_24;
wire q_21_25;
wire q_21_26;
wire q_21_27;
wire q_21_28;
wire q_21_29;
wire q_21_30;
wire q_21_31;
wire q_21_32;
wire q_21_33;
wire q_21_34;
wire q_21_35;
wire q_21_36;
wire q_21_37;
wire q_21_38;
wire q_21_39;
wire q_22_0;
wire q_22_1;
wire q_22_2;
wire q_22_3;
wire q_22_4;
wire q_22_5;
wire q_22_6;
wire q_22_7;
wire q_22_8;
wire q_22_9;
wire q_22_10;
wire q_22_11;
wire q_22_12;
wire q_22_13;
wire q_22_14;
wire q_22_15;
wire q_22_16;
wire q_22_17;
wire q_22_18;
wire q_22_19;
wire q_22_20;
wire q_22_21;
wire q_22_22;
wire q_22_23;
wire q_22_24;
wire q_22_25;
wire q_22_26;
wire q_22_27;
wire q_22_28;
wire q_22_29;
wire q_22_30;
wire q_22_31;
wire q_22_32;
wire q_22_33;
wire q_22_34;
wire q_22_35;
wire q_22_36;
wire q_22_37;
wire q_22_38;
wire q_22_39;
wire q_23_0;
wire q_23_1;
wire q_23_2;
wire q_23_3;
wire q_23_4;
wire q_23_5;
wire q_23_6;
wire q_23_7;
wire q_23_8;
wire q_23_9;
wire q_23_10;
wire q_23_11;
wire q_23_12;
wire q_23_13;
wire q_23_14;
wire q_23_15;
wire q_23_16;
wire q_23_17;
wire q_23_18;
wire q_23_19;
wire q_23_20;
wire q_23_21;
wire q_23_22;
wire q_23_23;
wire q_23_24;
wire q_23_25;
wire q_23_26;
wire q_23_27;
wire q_23_28;
wire q_23_29;
wire q_23_30;
wire q_23_31;
wire q_23_32;
wire q_23_33;
wire q_23_34;
wire q_23_35;
wire q_23_36;
wire q_23_37;
wire q_23_38;
wire q_23_39;
wire q_24_0;
wire q_24_1;
wire q_24_2;
wire q_24_3;
wire q_24_4;
wire q_24_5;
wire q_24_6;
wire q_24_7;
wire q_24_8;
wire q_24_9;
wire q_24_10;
wire q_24_11;
wire q_24_12;
wire q_24_13;
wire q_24_14;
wire q_24_15;
wire q_24_16;
wire q_24_17;
wire q_24_18;
wire q_24_19;
wire q_24_20;
wire q_24_21;
wire q_24_22;
wire q_24_23;
wire q_24_24;
wire q_24_25;
wire q_24_26;
wire q_24_27;
wire q_24_28;
wire q_24_29;
wire q_24_30;
wire q_24_31;
wire q_24_32;
wire q_24_33;
wire q_24_34;
wire q_24_35;
wire q_24_36;
wire q_24_37;
wire q_24_38;
wire q_24_39;
wire q_25_0;
wire q_25_1;
wire q_25_2;
wire q_25_3;
wire q_25_4;
wire q_25_5;
wire q_25_6;
wire q_25_7;
wire q_25_8;
wire q_25_9;
wire q_25_10;
wire q_25_11;
wire q_25_12;
wire q_25_13;
wire q_25_14;
wire q_25_15;
wire q_25_16;
wire q_25_17;
wire q_25_18;
wire q_25_19;
wire q_25_20;
wire q_25_21;
wire q_25_22;
wire q_25_23;
wire q_25_24;
wire q_25_25;
wire q_25_26;
wire q_25_27;
wire q_25_28;
wire q_25_29;
wire q_25_30;
wire q_25_31;
wire q_25_32;
wire q_25_33;
wire q_25_34;
wire q_25_35;
wire q_25_36;
wire q_25_37;
wire q_25_38;
wire q_25_39;
wire q_26_0;
wire q_26_1;
wire q_26_2;
wire q_26_3;
wire q_26_4;
wire q_26_5;
wire q_26_6;
wire q_26_7;
wire q_26_8;
wire q_26_9;
wire q_26_10;
wire q_26_11;
wire q_26_12;
wire q_26_13;
wire q_26_14;
wire q_26_15;
wire q_26_16;
wire q_26_17;
wire q_26_18;
wire q_26_19;
wire q_26_20;
wire q_26_21;
wire q_26_22;
wire q_26_23;
wire q_26_24;
wire q_26_25;
wire q_26_26;
wire q_26_27;
wire q_26_28;
wire q_26_29;
wire q_26_30;
wire q_26_31;
wire q_26_32;
wire q_26_33;
wire q_26_34;
wire q_26_35;
wire q_26_36;
wire q_26_37;
wire q_26_38;
wire q_26_39;
wire q_27_0;
wire q_27_1;
wire q_27_2;
wire q_27_3;
wire q_27_4;
wire q_27_5;
wire q_27_6;
wire q_27_7;
wire q_27_8;
wire q_27_9;
wire q_27_10;
wire q_27_11;
wire q_27_12;
wire q_27_13;
wire q_27_14;
wire q_27_15;
wire q_27_16;
wire q_27_17;
wire q_27_18;
wire q_27_19;
wire q_27_20;
wire q_27_21;
wire q_27_22;
wire q_27_23;
wire q_27_24;
wire q_27_25;
wire q_27_26;
wire q_27_27;
wire q_27_28;
wire q_27_29;
wire q_27_30;
wire q_27_31;
wire q_27_32;
wire q_27_33;
wire q_27_34;
wire q_27_35;
wire q_27_36;
wire q_27_37;
wire q_27_38;
wire q_27_39;
wire q_28_0;
wire q_28_1;
wire q_28_2;
wire q_28_3;
wire q_28_4;
wire q_28_5;
wire q_28_6;
wire q_28_7;
wire q_28_8;
wire q_28_9;
wire q_28_10;
wire q_28_11;
wire q_28_12;
wire q_28_13;
wire q_28_14;
wire q_28_15;
wire q_28_16;
wire q_28_17;
wire q_28_18;
wire q_28_19;
wire q_28_20;
wire q_28_21;
wire q_28_22;
wire q_28_23;
wire q_28_24;
wire q_28_25;
wire q_28_26;
wire q_28_27;
wire q_28_28;
wire q_28_29;
wire q_28_30;
wire q_28_31;
wire q_28_32;
wire q_28_33;
wire q_28_34;
wire q_28_35;
wire q_28_36;
wire q_28_37;
wire q_28_38;
wire q_28_39;
wire q_29_0;
wire q_29_1;
wire q_29_2;
wire q_29_3;
wire q_29_4;
wire q_29_5;
wire q_29_6;
wire q_29_7;
wire q_29_8;
wire q_29_9;
wire q_29_10;
wire q_29_11;
wire q_29_12;
wire q_29_13;
wire q_29_14;
wire q_29_15;
wire q_29_16;
wire q_29_17;
wire q_29_18;
wire q_29_19;
wire q_29_20;
wire q_29_21;
wire q_29_22;
wire q_29_23;
wire q_29_24;
wire q_29_25;
wire q_29_26;
wire q_29_27;
wire q_29_28;
wire q_29_29;
wire q_29_30;
wire q_29_31;
wire q_29_32;
wire q_29_33;
wire q_29_34;
wire q_29_35;
wire q_29_36;
wire q_29_37;
wire q_29_38;
wire q_29_39;
wire q_30_0;
wire q_30_1;
wire q_30_2;
wire q_30_3;
wire q_30_4;
wire q_30_5;
wire q_30_6;
wire q_30_7;
wire q_30_8;
wire q_30_9;
wire q_30_10;
wire q_30_11;
wire q_30_12;
wire q_30_13;
wire q_30_14;
wire q_30_15;
wire q_30_16;
wire q_30_17;
wire q_30_18;
wire q_30_19;
wire q_30_20;
wire q_30_21;
wire q_30_22;
wire q_30_23;
wire q_30_24;
wire q_30_25;
wire q_30_26;
wire q_30_27;
wire q_30_28;
wire q_30_29;
wire q_30_30;
wire q_30_31;
wire q_30_32;
wire q_30_33;
wire q_30_34;
wire q_30_35;
wire q_30_36;
wire q_30_37;
wire q_30_38;
wire q_30_39;
wire q_31_0;
wire q_31_1;
wire q_31_2;
wire q_31_3;
wire q_31_4;
wire q_31_5;
wire q_31_6;
wire q_31_7;
wire q_31_8;
wire q_31_9;
wire q_31_10;
wire q_31_11;
wire q_31_12;
wire q_31_13;
wire q_31_14;
wire q_31_15;
wire q_31_16;
wire q_31_17;
wire q_31_18;
wire q_31_19;
wire q_31_20;
wire q_31_21;
wire q_31_22;
wire q_31_23;
wire q_31_24;
wire q_31_25;
wire q_31_26;
wire q_31_27;
wire q_31_28;
wire q_31_29;
wire q_31_30;
wire q_31_31;
wire q_31_32;
wire q_31_33;
wire q_31_34;
wire q_31_35;
wire q_31_36;
wire q_31_37;
wire q_31_38;
wire q_31_39;
wire q_32_0;
wire q_32_1;
wire q_32_2;
wire q_32_3;
wire q_32_4;
wire q_32_5;
wire q_32_6;
wire q_32_7;
wire q_32_8;
wire q_32_9;
wire q_32_10;
wire q_32_11;
wire q_32_12;
wire q_32_13;
wire q_32_14;
wire q_32_15;
wire q_32_16;
wire q_32_17;
wire q_32_18;
wire q_32_19;
wire q_32_20;
wire q_32_21;
wire q_32_22;
wire q_32_23;
wire q_32_24;
wire q_32_25;
wire q_32_26;
wire q_32_27;
wire q_32_28;
wire q_32_29;
wire q_32_30;
wire q_32_31;
wire q_32_32;
wire q_32_33;
wire q_32_34;
wire q_32_35;
wire q_32_36;
wire q_32_37;
wire q_32_38;
wire q_32_39;
wire q_33_0;
wire q_33_1;
wire q_33_2;
wire q_33_3;
wire q_33_4;
wire q_33_5;
wire q_33_6;
wire q_33_7;
wire q_33_8;
wire q_33_9;
wire q_33_10;
wire q_33_11;
wire q_33_12;
wire q_33_13;
wire q_33_14;
wire q_33_15;
wire q_33_16;
wire q_33_17;
wire q_33_18;
wire q_33_19;
wire q_33_20;
wire q_33_21;
wire q_33_22;
wire q_33_23;
wire q_33_24;
wire q_33_25;
wire q_33_26;
wire q_33_27;
wire q_33_28;
wire q_33_29;
wire q_33_30;
wire q_33_31;
wire q_33_32;
wire q_33_33;
wire q_33_34;
wire q_33_35;
wire q_33_36;
wire q_33_37;
wire q_33_38;
wire q_33_39;
wire q_34_0;
wire q_34_1;
wire q_34_2;
wire q_34_3;
wire q_34_4;
wire q_34_5;
wire q_34_6;
wire q_34_7;
wire q_34_8;
wire q_34_9;
wire q_34_10;
wire q_34_11;
wire q_34_12;
wire q_34_13;
wire q_34_14;
wire q_34_15;
wire q_34_16;
wire q_34_17;
wire q_34_18;
wire q_34_19;
wire q_34_20;
wire q_34_21;
wire q_34_22;
wire q_34_23;
wire q_34_24;
wire q_34_25;
wire q_34_26;
wire q_34_27;
wire q_34_28;
wire q_34_29;
wire q_34_30;
wire q_34_31;
wire q_34_32;
wire q_34_33;
wire q_34_34;
wire q_34_35;
wire q_34_36;
wire q_34_37;
wire q_34_38;
wire q_34_39;
wire q_35_0;
wire q_35_1;
wire q_35_2;
wire q_35_3;
wire q_35_4;
wire q_35_5;
wire q_35_6;
wire q_35_7;
wire q_35_8;
wire q_35_9;
wire q_35_10;
wire q_35_11;
wire q_35_12;
wire q_35_13;
wire q_35_14;
wire q_35_15;
wire q_35_16;
wire q_35_17;
wire q_35_18;
wire q_35_19;
wire q_35_20;
wire q_35_21;
wire q_35_22;
wire q_35_23;
wire q_35_24;
wire q_35_25;
wire q_35_26;
wire q_35_27;
wire q_35_28;
wire q_35_29;
wire q_35_30;
wire q_35_31;
wire q_35_32;
wire q_35_33;
wire q_35_34;
wire q_35_35;
wire q_35_36;
wire q_35_37;
wire q_35_38;
wire q_35_39;
wire q_36_0;
wire q_36_1;
wire q_36_2;
wire q_36_3;
wire q_36_4;
wire q_36_5;
wire q_36_6;
wire q_36_7;
wire q_36_8;
wire q_36_9;
wire q_36_10;
wire q_36_11;
wire q_36_12;
wire q_36_13;
wire q_36_14;
wire q_36_15;
wire q_36_16;
wire q_36_17;
wire q_36_18;
wire q_36_19;
wire q_36_20;
wire q_36_21;
wire q_36_22;
wire q_36_23;
wire q_36_24;
wire q_36_25;
wire q_36_26;
wire q_36_27;
wire q_36_28;
wire q_36_29;
wire q_36_30;
wire q_36_31;
wire q_36_32;
wire q_36_33;
wire q_36_34;
wire q_36_35;
wire q_36_36;
wire q_36_37;
wire q_36_38;
wire q_36_39;
wire q_37_0;
wire q_37_1;
wire q_37_2;
wire q_37_3;
wire q_37_4;
wire q_37_5;
wire q_37_6;
wire q_37_7;
wire q_37_8;
wire q_37_9;
wire q_37_10;
wire q_37_11;
wire q_37_12;
wire q_37_13;
wire q_37_14;
wire q_37_15;
wire q_37_16;
wire q_37_17;
wire q_37_18;
wire q_37_19;
wire q_37_20;
wire q_37_21;
wire q_37_22;
wire q_37_23;
wire q_37_24;
wire q_37_25;
wire q_37_26;
wire q_37_27;
wire q_37_28;
wire q_37_29;
wire q_37_30;
wire q_37_31;
wire q_37_32;
wire q_37_33;
wire q_37_34;
wire q_37_35;
wire q_37_36;
wire q_37_37;
wire q_37_38;
wire q_37_39;
wire q_38_0;
wire q_38_1;
wire q_38_2;
wire q_38_3;
wire q_38_4;
wire q_38_5;
wire q_38_6;
wire q_38_7;
wire q_38_8;
wire q_38_9;
wire q_38_10;
wire q_38_11;
wire q_38_12;
wire q_38_13;
wire q_38_14;
wire q_38_15;
wire q_38_16;
wire q_38_17;
wire q_38_18;
wire q_38_19;
wire q_38_20;
wire q_38_21;
wire q_38_22;
wire q_38_23;
wire q_38_24;
wire q_38_25;
wire q_38_26;
wire q_38_27;
wire q_38_28;
wire q_38_29;
wire q_38_30;
wire q_38_31;
wire q_38_32;
wire q_38_33;
wire q_38_34;
wire q_38_35;
wire q_38_36;
wire q_38_37;
wire q_38_38;
wire q_38_39;
wire q_39_0;
wire q_39_1;
wire q_39_2;
wire q_39_3;
wire q_39_4;
wire q_39_5;
wire q_39_6;
wire q_39_7;
wire q_39_8;
wire q_39_9;
wire q_39_10;
wire q_39_11;
wire q_39_12;
wire q_39_13;
wire q_39_14;
wire q_39_15;
wire q_39_16;
wire q_39_17;
wire q_39_18;
wire q_39_19;
wire q_39_20;
wire q_39_21;
wire q_39_22;
wire q_39_23;
wire q_39_24;
wire q_39_25;
wire q_39_26;
wire q_39_27;
wire q_39_28;
wire q_39_29;
wire q_39_30;
wire q_39_31;
wire q_39_32;
wire q_39_33;
wire q_39_34;
wire q_39_35;
wire q_39_36;
wire q_39_37;
wire q_39_38;
wire q_39_39;

  wire q_0_minus1;
  assign q_0_minus1 = data_in[0];
  

  wire q_1_minus1;
  assign q_1_minus1 = data_in[1];
  

  wire q_2_minus1;
  assign q_2_minus1 = data_in[2];
  

  wire q_3_minus1;
  assign q_3_minus1 = data_in[3];
  

  wire q_4_minus1;
  assign q_4_minus1 = data_in[4];
  

  wire q_5_minus1;
  assign q_5_minus1 = data_in[5];
  

  wire q_6_minus1;
  assign q_6_minus1 = data_in[6];
  

  wire q_7_minus1;
  assign q_7_minus1 = data_in[7];
  

  wire q_8_minus1;
  assign q_8_minus1 = data_in[8];
  

  wire q_9_minus1;
  assign q_9_minus1 = data_in[9];
  

  wire q_10_minus1;
  assign q_10_minus1 = data_in[10];
  

  wire q_11_minus1;
  assign q_11_minus1 = data_in[11];
  

  wire q_12_minus1;
  assign q_12_minus1 = data_in[12];
  

  wire q_13_minus1;
  assign q_13_minus1 = data_in[13];
  

  wire q_14_minus1;
  assign q_14_minus1 = data_in[14];
  

  wire q_15_minus1;
  assign q_15_minus1 = data_in[15];
  

  wire q_16_minus1;
  assign q_16_minus1 = data_in[16];
  

  wire q_17_minus1;
  assign q_17_minus1 = data_in[17];
  

  wire q_18_minus1;
  assign q_18_minus1 = data_in[18];
  

  wire q_19_minus1;
  assign q_19_minus1 = data_in[19];
  

  wire q_20_minus1;
  assign q_20_minus1 = data_in[20];
  

  wire q_21_minus1;
  assign q_21_minus1 = data_in[21];
  

  wire q_22_minus1;
  assign q_22_minus1 = data_in[22];
  

  wire q_23_minus1;
  assign q_23_minus1 = data_in[23];
  

  wire q_24_minus1;
  assign q_24_minus1 = data_in[24];
  

  wire q_25_minus1;
  assign q_25_minus1 = data_in[25];
  

  wire q_26_minus1;
  assign q_26_minus1 = data_in[26];
  

  wire q_27_minus1;
  assign q_27_minus1 = data_in[27];
  

  wire q_28_minus1;
  assign q_28_minus1 = data_in[28];
  

  wire q_29_minus1;
  assign q_29_minus1 = data_in[29];
  

  wire q_30_minus1;
  assign q_30_minus1 = data_in[30];
  

  wire q_31_minus1;
  assign q_31_minus1 = data_in[31];
  

  wire q_32_minus1;
  assign q_32_minus1 = data_in[32];
  

  wire q_33_minus1;
  assign q_33_minus1 = data_in[33];
  

  wire q_34_minus1;
  assign q_34_minus1 = data_in[34];
  

  wire q_35_minus1;
  assign q_35_minus1 = data_in[35];
  

  wire q_36_minus1;
  assign q_36_minus1 = data_in[36];
  

  wire q_37_minus1;
  assign q_37_minus1 = data_in[37];
  

  wire q_38_minus1;
  assign q_38_minus1 = data_in[38];
  

  wire q_39_minus1;
  assign q_39_minus1 = data_in[39];
  

  assign data_out_internal[0] = q_39_0;
  

  assign data_out_internal[1] = q_39_1;
  

  assign data_out_internal[2] = q_39_2;
  

  assign data_out_internal[3] = q_39_3;
  

  assign data_out_internal[4] = q_39_4;
  

  assign data_out_internal[5] = q_39_5;
  

  assign data_out_internal[6] = q_39_6;
  

  assign data_out_internal[7] = q_39_7;
  

  assign data_out_internal[8] = q_39_8;
  

  assign data_out_internal[9] = q_39_9;
  

  assign data_out_internal[10] = q_39_10;
  

  assign data_out_internal[11] = q_39_11;
  

  assign data_out_internal[12] = q_39_12;
  

  assign data_out_internal[13] = q_39_13;
  

  assign data_out_internal[14] = q_39_14;
  

  assign data_out_internal[15] = q_39_15;
  

  assign data_out_internal[16] = q_39_16;
  

  assign data_out_internal[17] = q_39_17;
  

  assign data_out_internal[18] = q_39_18;
  

  assign data_out_internal[19] = q_39_19;
  

  assign data_out_internal[20] = q_39_20;
  

  assign data_out_internal[21] = q_39_21;
  

  assign data_out_internal[22] = q_39_22;
  

  assign data_out_internal[23] = q_39_23;
  

  assign data_out_internal[24] = q_39_24;
  

  assign data_out_internal[25] = q_39_25;
  

  assign data_out_internal[26] = q_39_26;
  

  assign data_out_internal[27] = q_39_27;
  

  assign data_out_internal[28] = q_39_28;
  

  assign data_out_internal[29] = q_39_29;
  

  assign data_out_internal[30] = q_39_30;
  

  assign data_out_internal[31] = q_39_31;
  

  assign data_out_internal[32] = q_39_32;
  

  assign data_out_internal[33] = q_39_33;
  

  assign data_out_internal[34] = q_39_34;
  

  assign data_out_internal[35] = q_39_35;
  

  assign data_out_internal[36] = q_39_36;
  

  assign data_out_internal[37] = q_39_37;
  

  assign data_out_internal[38] = q_39_38;
  

  assign data_out_internal[39] = q_39_39;
  

  wire q_minus1_0;
  assign q_minus1_0 = 1'b0;
  

  wire q_minus1_1;
  assign q_minus1_1 = 1'b0;
  

  wire q_minus1_2;
  assign q_minus1_2 = 1'b0;
  

  wire q_minus1_3;
  assign q_minus1_3 = 1'b0;
  

  wire q_minus1_4;
  assign q_minus1_4 = 1'b0;
  

  wire q_minus1_5;
  assign q_minus1_5 = 1'b0;
  

  wire q_minus1_6;
  assign q_minus1_6 = 1'b0;
  

  wire q_minus1_7;
  assign q_minus1_7 = 1'b0;
  

  wire q_minus1_8;
  assign q_minus1_8 = 1'b0;
  

  wire q_minus1_9;
  assign q_minus1_9 = 1'b0;
  

  wire q_minus1_10;
  assign q_minus1_10 = 1'b0;
  

  wire q_minus1_11;
  assign q_minus1_11 = 1'b0;
  

  wire q_minus1_12;
  assign q_minus1_12 = 1'b0;
  

  wire q_minus1_13;
  assign q_minus1_13 = 1'b0;
  

  wire q_minus1_14;
  assign q_minus1_14 = 1'b0;
  

  wire q_minus1_15;
  assign q_minus1_15 = 1'b0;
  

  wire q_minus1_16;
  assign q_minus1_16 = 1'b0;
  

  wire q_minus1_17;
  assign q_minus1_17 = 1'b0;
  

  wire q_minus1_18;
  assign q_minus1_18 = 1'b0;
  

  wire q_minus1_19;
  assign q_minus1_19 = 1'b0;
  

  wire q_minus1_20;
  assign q_minus1_20 = 1'b0;
  

  wire q_minus1_21;
  assign q_minus1_21 = 1'b0;
  

  wire q_minus1_22;
  assign q_minus1_22 = 1'b0;
  

  wire q_minus1_23;
  assign q_minus1_23 = 1'b0;
  

  wire q_minus1_24;
  assign q_minus1_24 = 1'b0;
  

  wire q_minus1_25;
  assign q_minus1_25 = 1'b0;
  

  wire q_minus1_26;
  assign q_minus1_26 = 1'b0;
  

  wire q_minus1_27;
  assign q_minus1_27 = 1'b0;
  

  wire q_minus1_28;
  assign q_minus1_28 = 1'b0;
  

  wire q_minus1_29;
  assign q_minus1_29 = 1'b0;
  

  wire q_minus1_30;
  assign q_minus1_30 = 1'b0;
  

  wire q_minus1_31;
  assign q_minus1_31 = 1'b0;
  

  wire q_minus1_32;
  assign q_minus1_32 = 1'b0;
  

  wire q_minus1_33;
  assign q_minus1_33 = 1'b0;
  

  wire q_minus1_34;
  assign q_minus1_34 = 1'b0;
  

  wire q_minus1_35;
  assign q_minus1_35 = 1'b0;
  

  wire q_minus1_36;
  assign q_minus1_36 = 1'b0;
  

  wire q_minus1_37;
  assign q_minus1_37 = 1'b0;
  

  wire q_minus1_38;
  assign q_minus1_38 = 1'b0;
  

  wire q_minus1_39;
  assign q_minus1_39 = 1'b0;
  

  flop_with_mux u_0_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_minus1),
    .d1(q_minus1_0),
    .q(q_0_0)
  );
  

  flop_with_mux u_0_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_0),
    .d1(q_minus1_1),
    .q(q_0_1)
  );
  

  flop_with_mux u_0_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_1),
    .d1(q_minus1_2),
    .q(q_0_2)
  );
  

  flop_with_mux u_0_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_2),
    .d1(q_minus1_3),
    .q(q_0_3)
  );
  

  flop_with_mux u_0_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_3),
    .d1(q_minus1_4),
    .q(q_0_4)
  );
  

  flop_with_mux u_0_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_4),
    .d1(q_minus1_5),
    .q(q_0_5)
  );
  

  flop_with_mux u_0_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_5),
    .d1(q_minus1_6),
    .q(q_0_6)
  );
  

  flop_with_mux u_0_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_6),
    .d1(q_minus1_7),
    .q(q_0_7)
  );
  

  flop_with_mux u_0_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_7),
    .d1(q_minus1_8),
    .q(q_0_8)
  );
  

  flop_with_mux u_0_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_8),
    .d1(q_minus1_9),
    .q(q_0_9)
  );
  

  flop_with_mux u_0_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_9),
    .d1(q_minus1_10),
    .q(q_0_10)
  );
  

  flop_with_mux u_0_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_10),
    .d1(q_minus1_11),
    .q(q_0_11)
  );
  

  flop_with_mux u_0_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_11),
    .d1(q_minus1_12),
    .q(q_0_12)
  );
  

  flop_with_mux u_0_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_12),
    .d1(q_minus1_13),
    .q(q_0_13)
  );
  

  flop_with_mux u_0_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_13),
    .d1(q_minus1_14),
    .q(q_0_14)
  );
  

  flop_with_mux u_0_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_14),
    .d1(q_minus1_15),
    .q(q_0_15)
  );
  

  flop_with_mux u_0_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_15),
    .d1(q_minus1_16),
    .q(q_0_16)
  );
  

  flop_with_mux u_0_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_16),
    .d1(q_minus1_17),
    .q(q_0_17)
  );
  

  flop_with_mux u_0_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_17),
    .d1(q_minus1_18),
    .q(q_0_18)
  );
  

  flop_with_mux u_0_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_18),
    .d1(q_minus1_19),
    .q(q_0_19)
  );
  

  flop_with_mux u_0_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_19),
    .d1(q_minus1_20),
    .q(q_0_20)
  );
  

  flop_with_mux u_0_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_20),
    .d1(q_minus1_21),
    .q(q_0_21)
  );
  

  flop_with_mux u_0_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_21),
    .d1(q_minus1_22),
    .q(q_0_22)
  );
  

  flop_with_mux u_0_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_22),
    .d1(q_minus1_23),
    .q(q_0_23)
  );
  

  flop_with_mux u_0_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_23),
    .d1(q_minus1_24),
    .q(q_0_24)
  );
  

  flop_with_mux u_0_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_24),
    .d1(q_minus1_25),
    .q(q_0_25)
  );
  

  flop_with_mux u_0_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_25),
    .d1(q_minus1_26),
    .q(q_0_26)
  );
  

  flop_with_mux u_0_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_26),
    .d1(q_minus1_27),
    .q(q_0_27)
  );
  

  flop_with_mux u_0_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_27),
    .d1(q_minus1_28),
    .q(q_0_28)
  );
  

  flop_with_mux u_0_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_28),
    .d1(q_minus1_29),
    .q(q_0_29)
  );
  

  flop_with_mux u_0_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_29),
    .d1(q_minus1_30),
    .q(q_0_30)
  );
  

  flop_with_mux u_0_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_30),
    .d1(q_minus1_31),
    .q(q_0_31)
  );
  

  flop_with_mux u_0_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_31),
    .d1(q_minus1_32),
    .q(q_0_32)
  );
  

  flop_with_mux u_0_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_32),
    .d1(q_minus1_33),
    .q(q_0_33)
  );
  

  flop_with_mux u_0_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_33),
    .d1(q_minus1_34),
    .q(q_0_34)
  );
  

  flop_with_mux u_0_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_34),
    .d1(q_minus1_35),
    .q(q_0_35)
  );
  

  flop_with_mux u_0_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_35),
    .d1(q_minus1_36),
    .q(q_0_36)
  );
  

  flop_with_mux u_0_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_36),
    .d1(q_minus1_37),
    .q(q_0_37)
  );
  

  flop_with_mux u_0_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_37),
    .d1(q_minus1_38),
    .q(q_0_38)
  );
  

  flop_with_mux u_0_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_0_38),
    .d1(q_minus1_39),
    .q(q_0_39)
  );
  

  flop_with_mux u_1_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_minus1),
    .d1(q_0_0),
    .q(q_1_0)
  );
  

  flop_with_mux u_1_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_0),
    .d1(q_0_1),
    .q(q_1_1)
  );
  

  flop_with_mux u_1_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_1),
    .d1(q_0_2),
    .q(q_1_2)
  );
  

  flop_with_mux u_1_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_2),
    .d1(q_0_3),
    .q(q_1_3)
  );
  

  flop_with_mux u_1_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_3),
    .d1(q_0_4),
    .q(q_1_4)
  );
  

  flop_with_mux u_1_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_4),
    .d1(q_0_5),
    .q(q_1_5)
  );
  

  flop_with_mux u_1_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_5),
    .d1(q_0_6),
    .q(q_1_6)
  );
  

  flop_with_mux u_1_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_6),
    .d1(q_0_7),
    .q(q_1_7)
  );
  

  flop_with_mux u_1_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_7),
    .d1(q_0_8),
    .q(q_1_8)
  );
  

  flop_with_mux u_1_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_8),
    .d1(q_0_9),
    .q(q_1_9)
  );
  

  flop_with_mux u_1_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_9),
    .d1(q_0_10),
    .q(q_1_10)
  );
  

  flop_with_mux u_1_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_10),
    .d1(q_0_11),
    .q(q_1_11)
  );
  

  flop_with_mux u_1_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_11),
    .d1(q_0_12),
    .q(q_1_12)
  );
  

  flop_with_mux u_1_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_12),
    .d1(q_0_13),
    .q(q_1_13)
  );
  

  flop_with_mux u_1_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_13),
    .d1(q_0_14),
    .q(q_1_14)
  );
  

  flop_with_mux u_1_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_14),
    .d1(q_0_15),
    .q(q_1_15)
  );
  

  flop_with_mux u_1_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_15),
    .d1(q_0_16),
    .q(q_1_16)
  );
  

  flop_with_mux u_1_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_16),
    .d1(q_0_17),
    .q(q_1_17)
  );
  

  flop_with_mux u_1_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_17),
    .d1(q_0_18),
    .q(q_1_18)
  );
  

  flop_with_mux u_1_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_18),
    .d1(q_0_19),
    .q(q_1_19)
  );
  

  flop_with_mux u_1_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_19),
    .d1(q_0_20),
    .q(q_1_20)
  );
  

  flop_with_mux u_1_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_20),
    .d1(q_0_21),
    .q(q_1_21)
  );
  

  flop_with_mux u_1_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_21),
    .d1(q_0_22),
    .q(q_1_22)
  );
  

  flop_with_mux u_1_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_22),
    .d1(q_0_23),
    .q(q_1_23)
  );
  

  flop_with_mux u_1_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_23),
    .d1(q_0_24),
    .q(q_1_24)
  );
  

  flop_with_mux u_1_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_24),
    .d1(q_0_25),
    .q(q_1_25)
  );
  

  flop_with_mux u_1_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_25),
    .d1(q_0_26),
    .q(q_1_26)
  );
  

  flop_with_mux u_1_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_26),
    .d1(q_0_27),
    .q(q_1_27)
  );
  

  flop_with_mux u_1_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_27),
    .d1(q_0_28),
    .q(q_1_28)
  );
  

  flop_with_mux u_1_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_28),
    .d1(q_0_29),
    .q(q_1_29)
  );
  

  flop_with_mux u_1_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_29),
    .d1(q_0_30),
    .q(q_1_30)
  );
  

  flop_with_mux u_1_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_30),
    .d1(q_0_31),
    .q(q_1_31)
  );
  

  flop_with_mux u_1_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_31),
    .d1(q_0_32),
    .q(q_1_32)
  );
  

  flop_with_mux u_1_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_32),
    .d1(q_0_33),
    .q(q_1_33)
  );
  

  flop_with_mux u_1_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_33),
    .d1(q_0_34),
    .q(q_1_34)
  );
  

  flop_with_mux u_1_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_34),
    .d1(q_0_35),
    .q(q_1_35)
  );
  

  flop_with_mux u_1_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_35),
    .d1(q_0_36),
    .q(q_1_36)
  );
  

  flop_with_mux u_1_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_36),
    .d1(q_0_37),
    .q(q_1_37)
  );
  

  flop_with_mux u_1_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_37),
    .d1(q_0_38),
    .q(q_1_38)
  );
  

  flop_with_mux u_1_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_1_38),
    .d1(q_0_39),
    .q(q_1_39)
  );
  

  flop_with_mux u_2_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_minus1),
    .d1(q_1_0),
    .q(q_2_0)
  );
  

  flop_with_mux u_2_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_0),
    .d1(q_1_1),
    .q(q_2_1)
  );
  

  flop_with_mux u_2_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_1),
    .d1(q_1_2),
    .q(q_2_2)
  );
  

  flop_with_mux u_2_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_2),
    .d1(q_1_3),
    .q(q_2_3)
  );
  

  flop_with_mux u_2_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_3),
    .d1(q_1_4),
    .q(q_2_4)
  );
  

  flop_with_mux u_2_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_4),
    .d1(q_1_5),
    .q(q_2_5)
  );
  

  flop_with_mux u_2_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_5),
    .d1(q_1_6),
    .q(q_2_6)
  );
  

  flop_with_mux u_2_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_6),
    .d1(q_1_7),
    .q(q_2_7)
  );
  

  flop_with_mux u_2_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_7),
    .d1(q_1_8),
    .q(q_2_8)
  );
  

  flop_with_mux u_2_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_8),
    .d1(q_1_9),
    .q(q_2_9)
  );
  

  flop_with_mux u_2_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_9),
    .d1(q_1_10),
    .q(q_2_10)
  );
  

  flop_with_mux u_2_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_10),
    .d1(q_1_11),
    .q(q_2_11)
  );
  

  flop_with_mux u_2_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_11),
    .d1(q_1_12),
    .q(q_2_12)
  );
  

  flop_with_mux u_2_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_12),
    .d1(q_1_13),
    .q(q_2_13)
  );
  

  flop_with_mux u_2_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_13),
    .d1(q_1_14),
    .q(q_2_14)
  );
  

  flop_with_mux u_2_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_14),
    .d1(q_1_15),
    .q(q_2_15)
  );
  

  flop_with_mux u_2_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_15),
    .d1(q_1_16),
    .q(q_2_16)
  );
  

  flop_with_mux u_2_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_16),
    .d1(q_1_17),
    .q(q_2_17)
  );
  

  flop_with_mux u_2_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_17),
    .d1(q_1_18),
    .q(q_2_18)
  );
  

  flop_with_mux u_2_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_18),
    .d1(q_1_19),
    .q(q_2_19)
  );
  

  flop_with_mux u_2_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_19),
    .d1(q_1_20),
    .q(q_2_20)
  );
  

  flop_with_mux u_2_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_20),
    .d1(q_1_21),
    .q(q_2_21)
  );
  

  flop_with_mux u_2_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_21),
    .d1(q_1_22),
    .q(q_2_22)
  );
  

  flop_with_mux u_2_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_22),
    .d1(q_1_23),
    .q(q_2_23)
  );
  

  flop_with_mux u_2_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_23),
    .d1(q_1_24),
    .q(q_2_24)
  );
  

  flop_with_mux u_2_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_24),
    .d1(q_1_25),
    .q(q_2_25)
  );
  

  flop_with_mux u_2_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_25),
    .d1(q_1_26),
    .q(q_2_26)
  );
  

  flop_with_mux u_2_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_26),
    .d1(q_1_27),
    .q(q_2_27)
  );
  

  flop_with_mux u_2_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_27),
    .d1(q_1_28),
    .q(q_2_28)
  );
  

  flop_with_mux u_2_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_28),
    .d1(q_1_29),
    .q(q_2_29)
  );
  

  flop_with_mux u_2_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_29),
    .d1(q_1_30),
    .q(q_2_30)
  );
  

  flop_with_mux u_2_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_30),
    .d1(q_1_31),
    .q(q_2_31)
  );
  

  flop_with_mux u_2_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_31),
    .d1(q_1_32),
    .q(q_2_32)
  );
  

  flop_with_mux u_2_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_32),
    .d1(q_1_33),
    .q(q_2_33)
  );
  

  flop_with_mux u_2_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_33),
    .d1(q_1_34),
    .q(q_2_34)
  );
  

  flop_with_mux u_2_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_34),
    .d1(q_1_35),
    .q(q_2_35)
  );
  

  flop_with_mux u_2_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_35),
    .d1(q_1_36),
    .q(q_2_36)
  );
  

  flop_with_mux u_2_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_36),
    .d1(q_1_37),
    .q(q_2_37)
  );
  

  flop_with_mux u_2_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_37),
    .d1(q_1_38),
    .q(q_2_38)
  );
  

  flop_with_mux u_2_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_2_38),
    .d1(q_1_39),
    .q(q_2_39)
  );
  

  flop_with_mux u_3_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_minus1),
    .d1(q_2_0),
    .q(q_3_0)
  );
  

  flop_with_mux u_3_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_0),
    .d1(q_2_1),
    .q(q_3_1)
  );
  

  flop_with_mux u_3_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_1),
    .d1(q_2_2),
    .q(q_3_2)
  );
  

  flop_with_mux u_3_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_2),
    .d1(q_2_3),
    .q(q_3_3)
  );
  

  flop_with_mux u_3_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_3),
    .d1(q_2_4),
    .q(q_3_4)
  );
  

  flop_with_mux u_3_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_4),
    .d1(q_2_5),
    .q(q_3_5)
  );
  

  flop_with_mux u_3_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_5),
    .d1(q_2_6),
    .q(q_3_6)
  );
  

  flop_with_mux u_3_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_6),
    .d1(q_2_7),
    .q(q_3_7)
  );
  

  flop_with_mux u_3_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_7),
    .d1(q_2_8),
    .q(q_3_8)
  );
  

  flop_with_mux u_3_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_8),
    .d1(q_2_9),
    .q(q_3_9)
  );
  

  flop_with_mux u_3_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_9),
    .d1(q_2_10),
    .q(q_3_10)
  );
  

  flop_with_mux u_3_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_10),
    .d1(q_2_11),
    .q(q_3_11)
  );
  

  flop_with_mux u_3_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_11),
    .d1(q_2_12),
    .q(q_3_12)
  );
  

  flop_with_mux u_3_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_12),
    .d1(q_2_13),
    .q(q_3_13)
  );
  

  flop_with_mux u_3_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_13),
    .d1(q_2_14),
    .q(q_3_14)
  );
  

  flop_with_mux u_3_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_14),
    .d1(q_2_15),
    .q(q_3_15)
  );
  

  flop_with_mux u_3_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_15),
    .d1(q_2_16),
    .q(q_3_16)
  );
  

  flop_with_mux u_3_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_16),
    .d1(q_2_17),
    .q(q_3_17)
  );
  

  flop_with_mux u_3_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_17),
    .d1(q_2_18),
    .q(q_3_18)
  );
  

  flop_with_mux u_3_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_18),
    .d1(q_2_19),
    .q(q_3_19)
  );
  

  flop_with_mux u_3_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_19),
    .d1(q_2_20),
    .q(q_3_20)
  );
  

  flop_with_mux u_3_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_20),
    .d1(q_2_21),
    .q(q_3_21)
  );
  

  flop_with_mux u_3_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_21),
    .d1(q_2_22),
    .q(q_3_22)
  );
  

  flop_with_mux u_3_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_22),
    .d1(q_2_23),
    .q(q_3_23)
  );
  

  flop_with_mux u_3_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_23),
    .d1(q_2_24),
    .q(q_3_24)
  );
  

  flop_with_mux u_3_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_24),
    .d1(q_2_25),
    .q(q_3_25)
  );
  

  flop_with_mux u_3_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_25),
    .d1(q_2_26),
    .q(q_3_26)
  );
  

  flop_with_mux u_3_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_26),
    .d1(q_2_27),
    .q(q_3_27)
  );
  

  flop_with_mux u_3_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_27),
    .d1(q_2_28),
    .q(q_3_28)
  );
  

  flop_with_mux u_3_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_28),
    .d1(q_2_29),
    .q(q_3_29)
  );
  

  flop_with_mux u_3_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_29),
    .d1(q_2_30),
    .q(q_3_30)
  );
  

  flop_with_mux u_3_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_30),
    .d1(q_2_31),
    .q(q_3_31)
  );
  

  flop_with_mux u_3_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_31),
    .d1(q_2_32),
    .q(q_3_32)
  );
  

  flop_with_mux u_3_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_32),
    .d1(q_2_33),
    .q(q_3_33)
  );
  

  flop_with_mux u_3_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_33),
    .d1(q_2_34),
    .q(q_3_34)
  );
  

  flop_with_mux u_3_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_34),
    .d1(q_2_35),
    .q(q_3_35)
  );
  

  flop_with_mux u_3_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_35),
    .d1(q_2_36),
    .q(q_3_36)
  );
  

  flop_with_mux u_3_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_36),
    .d1(q_2_37),
    .q(q_3_37)
  );
  

  flop_with_mux u_3_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_37),
    .d1(q_2_38),
    .q(q_3_38)
  );
  

  flop_with_mux u_3_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_3_38),
    .d1(q_2_39),
    .q(q_3_39)
  );
  

  flop_with_mux u_4_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_minus1),
    .d1(q_3_0),
    .q(q_4_0)
  );
  

  flop_with_mux u_4_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_0),
    .d1(q_3_1),
    .q(q_4_1)
  );
  

  flop_with_mux u_4_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_1),
    .d1(q_3_2),
    .q(q_4_2)
  );
  

  flop_with_mux u_4_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_2),
    .d1(q_3_3),
    .q(q_4_3)
  );
  

  flop_with_mux u_4_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_3),
    .d1(q_3_4),
    .q(q_4_4)
  );
  

  flop_with_mux u_4_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_4),
    .d1(q_3_5),
    .q(q_4_5)
  );
  

  flop_with_mux u_4_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_5),
    .d1(q_3_6),
    .q(q_4_6)
  );
  

  flop_with_mux u_4_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_6),
    .d1(q_3_7),
    .q(q_4_7)
  );
  

  flop_with_mux u_4_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_7),
    .d1(q_3_8),
    .q(q_4_8)
  );
  

  flop_with_mux u_4_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_8),
    .d1(q_3_9),
    .q(q_4_9)
  );
  

  flop_with_mux u_4_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_9),
    .d1(q_3_10),
    .q(q_4_10)
  );
  

  flop_with_mux u_4_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_10),
    .d1(q_3_11),
    .q(q_4_11)
  );
  

  flop_with_mux u_4_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_11),
    .d1(q_3_12),
    .q(q_4_12)
  );
  

  flop_with_mux u_4_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_12),
    .d1(q_3_13),
    .q(q_4_13)
  );
  

  flop_with_mux u_4_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_13),
    .d1(q_3_14),
    .q(q_4_14)
  );
  

  flop_with_mux u_4_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_14),
    .d1(q_3_15),
    .q(q_4_15)
  );
  

  flop_with_mux u_4_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_15),
    .d1(q_3_16),
    .q(q_4_16)
  );
  

  flop_with_mux u_4_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_16),
    .d1(q_3_17),
    .q(q_4_17)
  );
  

  flop_with_mux u_4_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_17),
    .d1(q_3_18),
    .q(q_4_18)
  );
  

  flop_with_mux u_4_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_18),
    .d1(q_3_19),
    .q(q_4_19)
  );
  

  flop_with_mux u_4_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_19),
    .d1(q_3_20),
    .q(q_4_20)
  );
  

  flop_with_mux u_4_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_20),
    .d1(q_3_21),
    .q(q_4_21)
  );
  

  flop_with_mux u_4_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_21),
    .d1(q_3_22),
    .q(q_4_22)
  );
  

  flop_with_mux u_4_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_22),
    .d1(q_3_23),
    .q(q_4_23)
  );
  

  flop_with_mux u_4_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_23),
    .d1(q_3_24),
    .q(q_4_24)
  );
  

  flop_with_mux u_4_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_24),
    .d1(q_3_25),
    .q(q_4_25)
  );
  

  flop_with_mux u_4_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_25),
    .d1(q_3_26),
    .q(q_4_26)
  );
  

  flop_with_mux u_4_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_26),
    .d1(q_3_27),
    .q(q_4_27)
  );
  

  flop_with_mux u_4_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_27),
    .d1(q_3_28),
    .q(q_4_28)
  );
  

  flop_with_mux u_4_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_28),
    .d1(q_3_29),
    .q(q_4_29)
  );
  

  flop_with_mux u_4_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_29),
    .d1(q_3_30),
    .q(q_4_30)
  );
  

  flop_with_mux u_4_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_30),
    .d1(q_3_31),
    .q(q_4_31)
  );
  

  flop_with_mux u_4_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_31),
    .d1(q_3_32),
    .q(q_4_32)
  );
  

  flop_with_mux u_4_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_32),
    .d1(q_3_33),
    .q(q_4_33)
  );
  

  flop_with_mux u_4_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_33),
    .d1(q_3_34),
    .q(q_4_34)
  );
  

  flop_with_mux u_4_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_34),
    .d1(q_3_35),
    .q(q_4_35)
  );
  

  flop_with_mux u_4_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_35),
    .d1(q_3_36),
    .q(q_4_36)
  );
  

  flop_with_mux u_4_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_36),
    .d1(q_3_37),
    .q(q_4_37)
  );
  

  flop_with_mux u_4_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_37),
    .d1(q_3_38),
    .q(q_4_38)
  );
  

  flop_with_mux u_4_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_4_38),
    .d1(q_3_39),
    .q(q_4_39)
  );
  

  flop_with_mux u_5_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_minus1),
    .d1(q_4_0),
    .q(q_5_0)
  );
  

  flop_with_mux u_5_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_0),
    .d1(q_4_1),
    .q(q_5_1)
  );
  

  flop_with_mux u_5_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_1),
    .d1(q_4_2),
    .q(q_5_2)
  );
  

  flop_with_mux u_5_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_2),
    .d1(q_4_3),
    .q(q_5_3)
  );
  

  flop_with_mux u_5_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_3),
    .d1(q_4_4),
    .q(q_5_4)
  );
  

  flop_with_mux u_5_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_4),
    .d1(q_4_5),
    .q(q_5_5)
  );
  

  flop_with_mux u_5_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_5),
    .d1(q_4_6),
    .q(q_5_6)
  );
  

  flop_with_mux u_5_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_6),
    .d1(q_4_7),
    .q(q_5_7)
  );
  

  flop_with_mux u_5_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_7),
    .d1(q_4_8),
    .q(q_5_8)
  );
  

  flop_with_mux u_5_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_8),
    .d1(q_4_9),
    .q(q_5_9)
  );
  

  flop_with_mux u_5_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_9),
    .d1(q_4_10),
    .q(q_5_10)
  );
  

  flop_with_mux u_5_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_10),
    .d1(q_4_11),
    .q(q_5_11)
  );
  

  flop_with_mux u_5_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_11),
    .d1(q_4_12),
    .q(q_5_12)
  );
  

  flop_with_mux u_5_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_12),
    .d1(q_4_13),
    .q(q_5_13)
  );
  

  flop_with_mux u_5_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_13),
    .d1(q_4_14),
    .q(q_5_14)
  );
  

  flop_with_mux u_5_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_14),
    .d1(q_4_15),
    .q(q_5_15)
  );
  

  flop_with_mux u_5_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_15),
    .d1(q_4_16),
    .q(q_5_16)
  );
  

  flop_with_mux u_5_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_16),
    .d1(q_4_17),
    .q(q_5_17)
  );
  

  flop_with_mux u_5_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_17),
    .d1(q_4_18),
    .q(q_5_18)
  );
  

  flop_with_mux u_5_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_18),
    .d1(q_4_19),
    .q(q_5_19)
  );
  

  flop_with_mux u_5_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_19),
    .d1(q_4_20),
    .q(q_5_20)
  );
  

  flop_with_mux u_5_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_20),
    .d1(q_4_21),
    .q(q_5_21)
  );
  

  flop_with_mux u_5_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_21),
    .d1(q_4_22),
    .q(q_5_22)
  );
  

  flop_with_mux u_5_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_22),
    .d1(q_4_23),
    .q(q_5_23)
  );
  

  flop_with_mux u_5_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_23),
    .d1(q_4_24),
    .q(q_5_24)
  );
  

  flop_with_mux u_5_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_24),
    .d1(q_4_25),
    .q(q_5_25)
  );
  

  flop_with_mux u_5_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_25),
    .d1(q_4_26),
    .q(q_5_26)
  );
  

  flop_with_mux u_5_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_26),
    .d1(q_4_27),
    .q(q_5_27)
  );
  

  flop_with_mux u_5_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_27),
    .d1(q_4_28),
    .q(q_5_28)
  );
  

  flop_with_mux u_5_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_28),
    .d1(q_4_29),
    .q(q_5_29)
  );
  

  flop_with_mux u_5_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_29),
    .d1(q_4_30),
    .q(q_5_30)
  );
  

  flop_with_mux u_5_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_30),
    .d1(q_4_31),
    .q(q_5_31)
  );
  

  flop_with_mux u_5_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_31),
    .d1(q_4_32),
    .q(q_5_32)
  );
  

  flop_with_mux u_5_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_32),
    .d1(q_4_33),
    .q(q_5_33)
  );
  

  flop_with_mux u_5_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_33),
    .d1(q_4_34),
    .q(q_5_34)
  );
  

  flop_with_mux u_5_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_34),
    .d1(q_4_35),
    .q(q_5_35)
  );
  

  flop_with_mux u_5_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_35),
    .d1(q_4_36),
    .q(q_5_36)
  );
  

  flop_with_mux u_5_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_36),
    .d1(q_4_37),
    .q(q_5_37)
  );
  

  flop_with_mux u_5_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_37),
    .d1(q_4_38),
    .q(q_5_38)
  );
  

  flop_with_mux u_5_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_5_38),
    .d1(q_4_39),
    .q(q_5_39)
  );
  

  flop_with_mux u_6_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_minus1),
    .d1(q_5_0),
    .q(q_6_0)
  );
  

  flop_with_mux u_6_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_0),
    .d1(q_5_1),
    .q(q_6_1)
  );
  

  flop_with_mux u_6_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_1),
    .d1(q_5_2),
    .q(q_6_2)
  );
  

  flop_with_mux u_6_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_2),
    .d1(q_5_3),
    .q(q_6_3)
  );
  

  flop_with_mux u_6_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_3),
    .d1(q_5_4),
    .q(q_6_4)
  );
  

  flop_with_mux u_6_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_4),
    .d1(q_5_5),
    .q(q_6_5)
  );
  

  flop_with_mux u_6_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_5),
    .d1(q_5_6),
    .q(q_6_6)
  );
  

  flop_with_mux u_6_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_6),
    .d1(q_5_7),
    .q(q_6_7)
  );
  

  flop_with_mux u_6_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_7),
    .d1(q_5_8),
    .q(q_6_8)
  );
  

  flop_with_mux u_6_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_8),
    .d1(q_5_9),
    .q(q_6_9)
  );
  

  flop_with_mux u_6_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_9),
    .d1(q_5_10),
    .q(q_6_10)
  );
  

  flop_with_mux u_6_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_10),
    .d1(q_5_11),
    .q(q_6_11)
  );
  

  flop_with_mux u_6_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_11),
    .d1(q_5_12),
    .q(q_6_12)
  );
  

  flop_with_mux u_6_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_12),
    .d1(q_5_13),
    .q(q_6_13)
  );
  

  flop_with_mux u_6_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_13),
    .d1(q_5_14),
    .q(q_6_14)
  );
  

  flop_with_mux u_6_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_14),
    .d1(q_5_15),
    .q(q_6_15)
  );
  

  flop_with_mux u_6_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_15),
    .d1(q_5_16),
    .q(q_6_16)
  );
  

  flop_with_mux u_6_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_16),
    .d1(q_5_17),
    .q(q_6_17)
  );
  

  flop_with_mux u_6_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_17),
    .d1(q_5_18),
    .q(q_6_18)
  );
  

  flop_with_mux u_6_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_18),
    .d1(q_5_19),
    .q(q_6_19)
  );
  

  flop_with_mux u_6_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_19),
    .d1(q_5_20),
    .q(q_6_20)
  );
  

  flop_with_mux u_6_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_20),
    .d1(q_5_21),
    .q(q_6_21)
  );
  

  flop_with_mux u_6_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_21),
    .d1(q_5_22),
    .q(q_6_22)
  );
  

  flop_with_mux u_6_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_22),
    .d1(q_5_23),
    .q(q_6_23)
  );
  

  flop_with_mux u_6_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_23),
    .d1(q_5_24),
    .q(q_6_24)
  );
  

  flop_with_mux u_6_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_24),
    .d1(q_5_25),
    .q(q_6_25)
  );
  

  flop_with_mux u_6_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_25),
    .d1(q_5_26),
    .q(q_6_26)
  );
  

  flop_with_mux u_6_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_26),
    .d1(q_5_27),
    .q(q_6_27)
  );
  

  flop_with_mux u_6_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_27),
    .d1(q_5_28),
    .q(q_6_28)
  );
  

  flop_with_mux u_6_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_28),
    .d1(q_5_29),
    .q(q_6_29)
  );
  

  flop_with_mux u_6_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_29),
    .d1(q_5_30),
    .q(q_6_30)
  );
  

  flop_with_mux u_6_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_30),
    .d1(q_5_31),
    .q(q_6_31)
  );
  

  flop_with_mux u_6_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_31),
    .d1(q_5_32),
    .q(q_6_32)
  );
  

  flop_with_mux u_6_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_32),
    .d1(q_5_33),
    .q(q_6_33)
  );
  

  flop_with_mux u_6_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_33),
    .d1(q_5_34),
    .q(q_6_34)
  );
  

  flop_with_mux u_6_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_34),
    .d1(q_5_35),
    .q(q_6_35)
  );
  

  flop_with_mux u_6_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_35),
    .d1(q_5_36),
    .q(q_6_36)
  );
  

  flop_with_mux u_6_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_36),
    .d1(q_5_37),
    .q(q_6_37)
  );
  

  flop_with_mux u_6_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_37),
    .d1(q_5_38),
    .q(q_6_38)
  );
  

  flop_with_mux u_6_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_6_38),
    .d1(q_5_39),
    .q(q_6_39)
  );
  

  flop_with_mux u_7_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_minus1),
    .d1(q_6_0),
    .q(q_7_0)
  );
  

  flop_with_mux u_7_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_0),
    .d1(q_6_1),
    .q(q_7_1)
  );
  

  flop_with_mux u_7_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_1),
    .d1(q_6_2),
    .q(q_7_2)
  );
  

  flop_with_mux u_7_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_2),
    .d1(q_6_3),
    .q(q_7_3)
  );
  

  flop_with_mux u_7_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_3),
    .d1(q_6_4),
    .q(q_7_4)
  );
  

  flop_with_mux u_7_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_4),
    .d1(q_6_5),
    .q(q_7_5)
  );
  

  flop_with_mux u_7_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_5),
    .d1(q_6_6),
    .q(q_7_6)
  );
  

  flop_with_mux u_7_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_6),
    .d1(q_6_7),
    .q(q_7_7)
  );
  

  flop_with_mux u_7_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_7),
    .d1(q_6_8),
    .q(q_7_8)
  );
  

  flop_with_mux u_7_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_8),
    .d1(q_6_9),
    .q(q_7_9)
  );
  

  flop_with_mux u_7_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_9),
    .d1(q_6_10),
    .q(q_7_10)
  );
  

  flop_with_mux u_7_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_10),
    .d1(q_6_11),
    .q(q_7_11)
  );
  

  flop_with_mux u_7_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_11),
    .d1(q_6_12),
    .q(q_7_12)
  );
  

  flop_with_mux u_7_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_12),
    .d1(q_6_13),
    .q(q_7_13)
  );
  

  flop_with_mux u_7_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_13),
    .d1(q_6_14),
    .q(q_7_14)
  );
  

  flop_with_mux u_7_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_14),
    .d1(q_6_15),
    .q(q_7_15)
  );
  

  flop_with_mux u_7_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_15),
    .d1(q_6_16),
    .q(q_7_16)
  );
  

  flop_with_mux u_7_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_16),
    .d1(q_6_17),
    .q(q_7_17)
  );
  

  flop_with_mux u_7_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_17),
    .d1(q_6_18),
    .q(q_7_18)
  );
  

  flop_with_mux u_7_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_18),
    .d1(q_6_19),
    .q(q_7_19)
  );
  

  flop_with_mux u_7_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_19),
    .d1(q_6_20),
    .q(q_7_20)
  );
  

  flop_with_mux u_7_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_20),
    .d1(q_6_21),
    .q(q_7_21)
  );
  

  flop_with_mux u_7_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_21),
    .d1(q_6_22),
    .q(q_7_22)
  );
  

  flop_with_mux u_7_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_22),
    .d1(q_6_23),
    .q(q_7_23)
  );
  

  flop_with_mux u_7_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_23),
    .d1(q_6_24),
    .q(q_7_24)
  );
  

  flop_with_mux u_7_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_24),
    .d1(q_6_25),
    .q(q_7_25)
  );
  

  flop_with_mux u_7_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_25),
    .d1(q_6_26),
    .q(q_7_26)
  );
  

  flop_with_mux u_7_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_26),
    .d1(q_6_27),
    .q(q_7_27)
  );
  

  flop_with_mux u_7_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_27),
    .d1(q_6_28),
    .q(q_7_28)
  );
  

  flop_with_mux u_7_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_28),
    .d1(q_6_29),
    .q(q_7_29)
  );
  

  flop_with_mux u_7_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_29),
    .d1(q_6_30),
    .q(q_7_30)
  );
  

  flop_with_mux u_7_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_30),
    .d1(q_6_31),
    .q(q_7_31)
  );
  

  flop_with_mux u_7_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_31),
    .d1(q_6_32),
    .q(q_7_32)
  );
  

  flop_with_mux u_7_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_32),
    .d1(q_6_33),
    .q(q_7_33)
  );
  

  flop_with_mux u_7_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_33),
    .d1(q_6_34),
    .q(q_7_34)
  );
  

  flop_with_mux u_7_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_34),
    .d1(q_6_35),
    .q(q_7_35)
  );
  

  flop_with_mux u_7_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_35),
    .d1(q_6_36),
    .q(q_7_36)
  );
  

  flop_with_mux u_7_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_36),
    .d1(q_6_37),
    .q(q_7_37)
  );
  

  flop_with_mux u_7_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_37),
    .d1(q_6_38),
    .q(q_7_38)
  );
  

  flop_with_mux u_7_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_7_38),
    .d1(q_6_39),
    .q(q_7_39)
  );
  

  flop_with_mux u_8_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_minus1),
    .d1(q_7_0),
    .q(q_8_0)
  );
  

  flop_with_mux u_8_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_0),
    .d1(q_7_1),
    .q(q_8_1)
  );
  

  flop_with_mux u_8_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_1),
    .d1(q_7_2),
    .q(q_8_2)
  );
  

  flop_with_mux u_8_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_2),
    .d1(q_7_3),
    .q(q_8_3)
  );
  

  flop_with_mux u_8_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_3),
    .d1(q_7_4),
    .q(q_8_4)
  );
  

  flop_with_mux u_8_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_4),
    .d1(q_7_5),
    .q(q_8_5)
  );
  

  flop_with_mux u_8_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_5),
    .d1(q_7_6),
    .q(q_8_6)
  );
  

  flop_with_mux u_8_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_6),
    .d1(q_7_7),
    .q(q_8_7)
  );
  

  flop_with_mux u_8_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_7),
    .d1(q_7_8),
    .q(q_8_8)
  );
  

  flop_with_mux u_8_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_8),
    .d1(q_7_9),
    .q(q_8_9)
  );
  

  flop_with_mux u_8_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_9),
    .d1(q_7_10),
    .q(q_8_10)
  );
  

  flop_with_mux u_8_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_10),
    .d1(q_7_11),
    .q(q_8_11)
  );
  

  flop_with_mux u_8_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_11),
    .d1(q_7_12),
    .q(q_8_12)
  );
  

  flop_with_mux u_8_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_12),
    .d1(q_7_13),
    .q(q_8_13)
  );
  

  flop_with_mux u_8_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_13),
    .d1(q_7_14),
    .q(q_8_14)
  );
  

  flop_with_mux u_8_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_14),
    .d1(q_7_15),
    .q(q_8_15)
  );
  

  flop_with_mux u_8_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_15),
    .d1(q_7_16),
    .q(q_8_16)
  );
  

  flop_with_mux u_8_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_16),
    .d1(q_7_17),
    .q(q_8_17)
  );
  

  flop_with_mux u_8_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_17),
    .d1(q_7_18),
    .q(q_8_18)
  );
  

  flop_with_mux u_8_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_18),
    .d1(q_7_19),
    .q(q_8_19)
  );
  

  flop_with_mux u_8_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_19),
    .d1(q_7_20),
    .q(q_8_20)
  );
  

  flop_with_mux u_8_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_20),
    .d1(q_7_21),
    .q(q_8_21)
  );
  

  flop_with_mux u_8_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_21),
    .d1(q_7_22),
    .q(q_8_22)
  );
  

  flop_with_mux u_8_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_22),
    .d1(q_7_23),
    .q(q_8_23)
  );
  

  flop_with_mux u_8_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_23),
    .d1(q_7_24),
    .q(q_8_24)
  );
  

  flop_with_mux u_8_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_24),
    .d1(q_7_25),
    .q(q_8_25)
  );
  

  flop_with_mux u_8_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_25),
    .d1(q_7_26),
    .q(q_8_26)
  );
  

  flop_with_mux u_8_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_26),
    .d1(q_7_27),
    .q(q_8_27)
  );
  

  flop_with_mux u_8_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_27),
    .d1(q_7_28),
    .q(q_8_28)
  );
  

  flop_with_mux u_8_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_28),
    .d1(q_7_29),
    .q(q_8_29)
  );
  

  flop_with_mux u_8_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_29),
    .d1(q_7_30),
    .q(q_8_30)
  );
  

  flop_with_mux u_8_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_30),
    .d1(q_7_31),
    .q(q_8_31)
  );
  

  flop_with_mux u_8_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_31),
    .d1(q_7_32),
    .q(q_8_32)
  );
  

  flop_with_mux u_8_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_32),
    .d1(q_7_33),
    .q(q_8_33)
  );
  

  flop_with_mux u_8_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_33),
    .d1(q_7_34),
    .q(q_8_34)
  );
  

  flop_with_mux u_8_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_34),
    .d1(q_7_35),
    .q(q_8_35)
  );
  

  flop_with_mux u_8_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_35),
    .d1(q_7_36),
    .q(q_8_36)
  );
  

  flop_with_mux u_8_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_36),
    .d1(q_7_37),
    .q(q_8_37)
  );
  

  flop_with_mux u_8_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_37),
    .d1(q_7_38),
    .q(q_8_38)
  );
  

  flop_with_mux u_8_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_8_38),
    .d1(q_7_39),
    .q(q_8_39)
  );
  

  flop_with_mux u_9_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_minus1),
    .d1(q_8_0),
    .q(q_9_0)
  );
  

  flop_with_mux u_9_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_0),
    .d1(q_8_1),
    .q(q_9_1)
  );
  

  flop_with_mux u_9_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_1),
    .d1(q_8_2),
    .q(q_9_2)
  );
  

  flop_with_mux u_9_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_2),
    .d1(q_8_3),
    .q(q_9_3)
  );
  

  flop_with_mux u_9_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_3),
    .d1(q_8_4),
    .q(q_9_4)
  );
  

  flop_with_mux u_9_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_4),
    .d1(q_8_5),
    .q(q_9_5)
  );
  

  flop_with_mux u_9_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_5),
    .d1(q_8_6),
    .q(q_9_6)
  );
  

  flop_with_mux u_9_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_6),
    .d1(q_8_7),
    .q(q_9_7)
  );
  

  flop_with_mux u_9_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_7),
    .d1(q_8_8),
    .q(q_9_8)
  );
  

  flop_with_mux u_9_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_8),
    .d1(q_8_9),
    .q(q_9_9)
  );
  

  flop_with_mux u_9_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_9),
    .d1(q_8_10),
    .q(q_9_10)
  );
  

  flop_with_mux u_9_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_10),
    .d1(q_8_11),
    .q(q_9_11)
  );
  

  flop_with_mux u_9_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_11),
    .d1(q_8_12),
    .q(q_9_12)
  );
  

  flop_with_mux u_9_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_12),
    .d1(q_8_13),
    .q(q_9_13)
  );
  

  flop_with_mux u_9_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_13),
    .d1(q_8_14),
    .q(q_9_14)
  );
  

  flop_with_mux u_9_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_14),
    .d1(q_8_15),
    .q(q_9_15)
  );
  

  flop_with_mux u_9_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_15),
    .d1(q_8_16),
    .q(q_9_16)
  );
  

  flop_with_mux u_9_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_16),
    .d1(q_8_17),
    .q(q_9_17)
  );
  

  flop_with_mux u_9_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_17),
    .d1(q_8_18),
    .q(q_9_18)
  );
  

  flop_with_mux u_9_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_18),
    .d1(q_8_19),
    .q(q_9_19)
  );
  

  flop_with_mux u_9_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_19),
    .d1(q_8_20),
    .q(q_9_20)
  );
  

  flop_with_mux u_9_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_20),
    .d1(q_8_21),
    .q(q_9_21)
  );
  

  flop_with_mux u_9_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_21),
    .d1(q_8_22),
    .q(q_9_22)
  );
  

  flop_with_mux u_9_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_22),
    .d1(q_8_23),
    .q(q_9_23)
  );
  

  flop_with_mux u_9_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_23),
    .d1(q_8_24),
    .q(q_9_24)
  );
  

  flop_with_mux u_9_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_24),
    .d1(q_8_25),
    .q(q_9_25)
  );
  

  flop_with_mux u_9_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_25),
    .d1(q_8_26),
    .q(q_9_26)
  );
  

  flop_with_mux u_9_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_26),
    .d1(q_8_27),
    .q(q_9_27)
  );
  

  flop_with_mux u_9_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_27),
    .d1(q_8_28),
    .q(q_9_28)
  );
  

  flop_with_mux u_9_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_28),
    .d1(q_8_29),
    .q(q_9_29)
  );
  

  flop_with_mux u_9_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_29),
    .d1(q_8_30),
    .q(q_9_30)
  );
  

  flop_with_mux u_9_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_30),
    .d1(q_8_31),
    .q(q_9_31)
  );
  

  flop_with_mux u_9_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_31),
    .d1(q_8_32),
    .q(q_9_32)
  );
  

  flop_with_mux u_9_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_32),
    .d1(q_8_33),
    .q(q_9_33)
  );
  

  flop_with_mux u_9_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_33),
    .d1(q_8_34),
    .q(q_9_34)
  );
  

  flop_with_mux u_9_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_34),
    .d1(q_8_35),
    .q(q_9_35)
  );
  

  flop_with_mux u_9_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_35),
    .d1(q_8_36),
    .q(q_9_36)
  );
  

  flop_with_mux u_9_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_36),
    .d1(q_8_37),
    .q(q_9_37)
  );
  

  flop_with_mux u_9_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_37),
    .d1(q_8_38),
    .q(q_9_38)
  );
  

  flop_with_mux u_9_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_9_38),
    .d1(q_8_39),
    .q(q_9_39)
  );
  

  flop_with_mux u_10_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_minus1),
    .d1(q_9_0),
    .q(q_10_0)
  );
  

  flop_with_mux u_10_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_0),
    .d1(q_9_1),
    .q(q_10_1)
  );
  

  flop_with_mux u_10_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_1),
    .d1(q_9_2),
    .q(q_10_2)
  );
  

  flop_with_mux u_10_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_2),
    .d1(q_9_3),
    .q(q_10_3)
  );
  

  flop_with_mux u_10_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_3),
    .d1(q_9_4),
    .q(q_10_4)
  );
  

  flop_with_mux u_10_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_4),
    .d1(q_9_5),
    .q(q_10_5)
  );
  

  flop_with_mux u_10_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_5),
    .d1(q_9_6),
    .q(q_10_6)
  );
  

  flop_with_mux u_10_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_6),
    .d1(q_9_7),
    .q(q_10_7)
  );
  

  flop_with_mux u_10_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_7),
    .d1(q_9_8),
    .q(q_10_8)
  );
  

  flop_with_mux u_10_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_8),
    .d1(q_9_9),
    .q(q_10_9)
  );
  

  flop_with_mux u_10_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_9),
    .d1(q_9_10),
    .q(q_10_10)
  );
  

  flop_with_mux u_10_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_10),
    .d1(q_9_11),
    .q(q_10_11)
  );
  

  flop_with_mux u_10_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_11),
    .d1(q_9_12),
    .q(q_10_12)
  );
  

  flop_with_mux u_10_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_12),
    .d1(q_9_13),
    .q(q_10_13)
  );
  

  flop_with_mux u_10_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_13),
    .d1(q_9_14),
    .q(q_10_14)
  );
  

  flop_with_mux u_10_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_14),
    .d1(q_9_15),
    .q(q_10_15)
  );
  

  flop_with_mux u_10_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_15),
    .d1(q_9_16),
    .q(q_10_16)
  );
  

  flop_with_mux u_10_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_16),
    .d1(q_9_17),
    .q(q_10_17)
  );
  

  flop_with_mux u_10_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_17),
    .d1(q_9_18),
    .q(q_10_18)
  );
  

  flop_with_mux u_10_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_18),
    .d1(q_9_19),
    .q(q_10_19)
  );
  

  flop_with_mux u_10_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_19),
    .d1(q_9_20),
    .q(q_10_20)
  );
  

  flop_with_mux u_10_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_20),
    .d1(q_9_21),
    .q(q_10_21)
  );
  

  flop_with_mux u_10_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_21),
    .d1(q_9_22),
    .q(q_10_22)
  );
  

  flop_with_mux u_10_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_22),
    .d1(q_9_23),
    .q(q_10_23)
  );
  

  flop_with_mux u_10_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_23),
    .d1(q_9_24),
    .q(q_10_24)
  );
  

  flop_with_mux u_10_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_24),
    .d1(q_9_25),
    .q(q_10_25)
  );
  

  flop_with_mux u_10_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_25),
    .d1(q_9_26),
    .q(q_10_26)
  );
  

  flop_with_mux u_10_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_26),
    .d1(q_9_27),
    .q(q_10_27)
  );
  

  flop_with_mux u_10_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_27),
    .d1(q_9_28),
    .q(q_10_28)
  );
  

  flop_with_mux u_10_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_28),
    .d1(q_9_29),
    .q(q_10_29)
  );
  

  flop_with_mux u_10_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_29),
    .d1(q_9_30),
    .q(q_10_30)
  );
  

  flop_with_mux u_10_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_30),
    .d1(q_9_31),
    .q(q_10_31)
  );
  

  flop_with_mux u_10_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_31),
    .d1(q_9_32),
    .q(q_10_32)
  );
  

  flop_with_mux u_10_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_32),
    .d1(q_9_33),
    .q(q_10_33)
  );
  

  flop_with_mux u_10_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_33),
    .d1(q_9_34),
    .q(q_10_34)
  );
  

  flop_with_mux u_10_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_34),
    .d1(q_9_35),
    .q(q_10_35)
  );
  

  flop_with_mux u_10_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_35),
    .d1(q_9_36),
    .q(q_10_36)
  );
  

  flop_with_mux u_10_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_36),
    .d1(q_9_37),
    .q(q_10_37)
  );
  

  flop_with_mux u_10_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_37),
    .d1(q_9_38),
    .q(q_10_38)
  );
  

  flop_with_mux u_10_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_10_38),
    .d1(q_9_39),
    .q(q_10_39)
  );
  

  flop_with_mux u_11_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_minus1),
    .d1(q_10_0),
    .q(q_11_0)
  );
  

  flop_with_mux u_11_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_0),
    .d1(q_10_1),
    .q(q_11_1)
  );
  

  flop_with_mux u_11_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_1),
    .d1(q_10_2),
    .q(q_11_2)
  );
  

  flop_with_mux u_11_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_2),
    .d1(q_10_3),
    .q(q_11_3)
  );
  

  flop_with_mux u_11_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_3),
    .d1(q_10_4),
    .q(q_11_4)
  );
  

  flop_with_mux u_11_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_4),
    .d1(q_10_5),
    .q(q_11_5)
  );
  

  flop_with_mux u_11_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_5),
    .d1(q_10_6),
    .q(q_11_6)
  );
  

  flop_with_mux u_11_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_6),
    .d1(q_10_7),
    .q(q_11_7)
  );
  

  flop_with_mux u_11_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_7),
    .d1(q_10_8),
    .q(q_11_8)
  );
  

  flop_with_mux u_11_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_8),
    .d1(q_10_9),
    .q(q_11_9)
  );
  

  flop_with_mux u_11_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_9),
    .d1(q_10_10),
    .q(q_11_10)
  );
  

  flop_with_mux u_11_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_10),
    .d1(q_10_11),
    .q(q_11_11)
  );
  

  flop_with_mux u_11_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_11),
    .d1(q_10_12),
    .q(q_11_12)
  );
  

  flop_with_mux u_11_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_12),
    .d1(q_10_13),
    .q(q_11_13)
  );
  

  flop_with_mux u_11_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_13),
    .d1(q_10_14),
    .q(q_11_14)
  );
  

  flop_with_mux u_11_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_14),
    .d1(q_10_15),
    .q(q_11_15)
  );
  

  flop_with_mux u_11_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_15),
    .d1(q_10_16),
    .q(q_11_16)
  );
  

  flop_with_mux u_11_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_16),
    .d1(q_10_17),
    .q(q_11_17)
  );
  

  flop_with_mux u_11_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_17),
    .d1(q_10_18),
    .q(q_11_18)
  );
  

  flop_with_mux u_11_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_18),
    .d1(q_10_19),
    .q(q_11_19)
  );
  

  flop_with_mux u_11_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_19),
    .d1(q_10_20),
    .q(q_11_20)
  );
  

  flop_with_mux u_11_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_20),
    .d1(q_10_21),
    .q(q_11_21)
  );
  

  flop_with_mux u_11_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_21),
    .d1(q_10_22),
    .q(q_11_22)
  );
  

  flop_with_mux u_11_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_22),
    .d1(q_10_23),
    .q(q_11_23)
  );
  

  flop_with_mux u_11_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_23),
    .d1(q_10_24),
    .q(q_11_24)
  );
  

  flop_with_mux u_11_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_24),
    .d1(q_10_25),
    .q(q_11_25)
  );
  

  flop_with_mux u_11_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_25),
    .d1(q_10_26),
    .q(q_11_26)
  );
  

  flop_with_mux u_11_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_26),
    .d1(q_10_27),
    .q(q_11_27)
  );
  

  flop_with_mux u_11_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_27),
    .d1(q_10_28),
    .q(q_11_28)
  );
  

  flop_with_mux u_11_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_28),
    .d1(q_10_29),
    .q(q_11_29)
  );
  

  flop_with_mux u_11_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_29),
    .d1(q_10_30),
    .q(q_11_30)
  );
  

  flop_with_mux u_11_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_30),
    .d1(q_10_31),
    .q(q_11_31)
  );
  

  flop_with_mux u_11_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_31),
    .d1(q_10_32),
    .q(q_11_32)
  );
  

  flop_with_mux u_11_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_32),
    .d1(q_10_33),
    .q(q_11_33)
  );
  

  flop_with_mux u_11_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_33),
    .d1(q_10_34),
    .q(q_11_34)
  );
  

  flop_with_mux u_11_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_34),
    .d1(q_10_35),
    .q(q_11_35)
  );
  

  flop_with_mux u_11_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_35),
    .d1(q_10_36),
    .q(q_11_36)
  );
  

  flop_with_mux u_11_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_36),
    .d1(q_10_37),
    .q(q_11_37)
  );
  

  flop_with_mux u_11_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_37),
    .d1(q_10_38),
    .q(q_11_38)
  );
  

  flop_with_mux u_11_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_11_38),
    .d1(q_10_39),
    .q(q_11_39)
  );
  

  flop_with_mux u_12_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_minus1),
    .d1(q_11_0),
    .q(q_12_0)
  );
  

  flop_with_mux u_12_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_0),
    .d1(q_11_1),
    .q(q_12_1)
  );
  

  flop_with_mux u_12_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_1),
    .d1(q_11_2),
    .q(q_12_2)
  );
  

  flop_with_mux u_12_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_2),
    .d1(q_11_3),
    .q(q_12_3)
  );
  

  flop_with_mux u_12_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_3),
    .d1(q_11_4),
    .q(q_12_4)
  );
  

  flop_with_mux u_12_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_4),
    .d1(q_11_5),
    .q(q_12_5)
  );
  

  flop_with_mux u_12_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_5),
    .d1(q_11_6),
    .q(q_12_6)
  );
  

  flop_with_mux u_12_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_6),
    .d1(q_11_7),
    .q(q_12_7)
  );
  

  flop_with_mux u_12_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_7),
    .d1(q_11_8),
    .q(q_12_8)
  );
  

  flop_with_mux u_12_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_8),
    .d1(q_11_9),
    .q(q_12_9)
  );
  

  flop_with_mux u_12_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_9),
    .d1(q_11_10),
    .q(q_12_10)
  );
  

  flop_with_mux u_12_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_10),
    .d1(q_11_11),
    .q(q_12_11)
  );
  

  flop_with_mux u_12_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_11),
    .d1(q_11_12),
    .q(q_12_12)
  );
  

  flop_with_mux u_12_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_12),
    .d1(q_11_13),
    .q(q_12_13)
  );
  

  flop_with_mux u_12_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_13),
    .d1(q_11_14),
    .q(q_12_14)
  );
  

  flop_with_mux u_12_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_14),
    .d1(q_11_15),
    .q(q_12_15)
  );
  

  flop_with_mux u_12_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_15),
    .d1(q_11_16),
    .q(q_12_16)
  );
  

  flop_with_mux u_12_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_16),
    .d1(q_11_17),
    .q(q_12_17)
  );
  

  flop_with_mux u_12_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_17),
    .d1(q_11_18),
    .q(q_12_18)
  );
  

  flop_with_mux u_12_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_18),
    .d1(q_11_19),
    .q(q_12_19)
  );
  

  flop_with_mux u_12_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_19),
    .d1(q_11_20),
    .q(q_12_20)
  );
  

  flop_with_mux u_12_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_20),
    .d1(q_11_21),
    .q(q_12_21)
  );
  

  flop_with_mux u_12_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_21),
    .d1(q_11_22),
    .q(q_12_22)
  );
  

  flop_with_mux u_12_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_22),
    .d1(q_11_23),
    .q(q_12_23)
  );
  

  flop_with_mux u_12_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_23),
    .d1(q_11_24),
    .q(q_12_24)
  );
  

  flop_with_mux u_12_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_24),
    .d1(q_11_25),
    .q(q_12_25)
  );
  

  flop_with_mux u_12_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_25),
    .d1(q_11_26),
    .q(q_12_26)
  );
  

  flop_with_mux u_12_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_26),
    .d1(q_11_27),
    .q(q_12_27)
  );
  

  flop_with_mux u_12_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_27),
    .d1(q_11_28),
    .q(q_12_28)
  );
  

  flop_with_mux u_12_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_28),
    .d1(q_11_29),
    .q(q_12_29)
  );
  

  flop_with_mux u_12_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_29),
    .d1(q_11_30),
    .q(q_12_30)
  );
  

  flop_with_mux u_12_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_30),
    .d1(q_11_31),
    .q(q_12_31)
  );
  

  flop_with_mux u_12_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_31),
    .d1(q_11_32),
    .q(q_12_32)
  );
  

  flop_with_mux u_12_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_32),
    .d1(q_11_33),
    .q(q_12_33)
  );
  

  flop_with_mux u_12_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_33),
    .d1(q_11_34),
    .q(q_12_34)
  );
  

  flop_with_mux u_12_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_34),
    .d1(q_11_35),
    .q(q_12_35)
  );
  

  flop_with_mux u_12_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_35),
    .d1(q_11_36),
    .q(q_12_36)
  );
  

  flop_with_mux u_12_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_36),
    .d1(q_11_37),
    .q(q_12_37)
  );
  

  flop_with_mux u_12_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_37),
    .d1(q_11_38),
    .q(q_12_38)
  );
  

  flop_with_mux u_12_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_12_38),
    .d1(q_11_39),
    .q(q_12_39)
  );
  

  flop_with_mux u_13_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_minus1),
    .d1(q_12_0),
    .q(q_13_0)
  );
  

  flop_with_mux u_13_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_0),
    .d1(q_12_1),
    .q(q_13_1)
  );
  

  flop_with_mux u_13_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_1),
    .d1(q_12_2),
    .q(q_13_2)
  );
  

  flop_with_mux u_13_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_2),
    .d1(q_12_3),
    .q(q_13_3)
  );
  

  flop_with_mux u_13_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_3),
    .d1(q_12_4),
    .q(q_13_4)
  );
  

  flop_with_mux u_13_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_4),
    .d1(q_12_5),
    .q(q_13_5)
  );
  

  flop_with_mux u_13_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_5),
    .d1(q_12_6),
    .q(q_13_6)
  );
  

  flop_with_mux u_13_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_6),
    .d1(q_12_7),
    .q(q_13_7)
  );
  

  flop_with_mux u_13_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_7),
    .d1(q_12_8),
    .q(q_13_8)
  );
  

  flop_with_mux u_13_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_8),
    .d1(q_12_9),
    .q(q_13_9)
  );
  

  flop_with_mux u_13_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_9),
    .d1(q_12_10),
    .q(q_13_10)
  );
  

  flop_with_mux u_13_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_10),
    .d1(q_12_11),
    .q(q_13_11)
  );
  

  flop_with_mux u_13_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_11),
    .d1(q_12_12),
    .q(q_13_12)
  );
  

  flop_with_mux u_13_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_12),
    .d1(q_12_13),
    .q(q_13_13)
  );
  

  flop_with_mux u_13_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_13),
    .d1(q_12_14),
    .q(q_13_14)
  );
  

  flop_with_mux u_13_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_14),
    .d1(q_12_15),
    .q(q_13_15)
  );
  

  flop_with_mux u_13_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_15),
    .d1(q_12_16),
    .q(q_13_16)
  );
  

  flop_with_mux u_13_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_16),
    .d1(q_12_17),
    .q(q_13_17)
  );
  

  flop_with_mux u_13_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_17),
    .d1(q_12_18),
    .q(q_13_18)
  );
  

  flop_with_mux u_13_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_18),
    .d1(q_12_19),
    .q(q_13_19)
  );
  

  flop_with_mux u_13_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_19),
    .d1(q_12_20),
    .q(q_13_20)
  );
  

  flop_with_mux u_13_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_20),
    .d1(q_12_21),
    .q(q_13_21)
  );
  

  flop_with_mux u_13_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_21),
    .d1(q_12_22),
    .q(q_13_22)
  );
  

  flop_with_mux u_13_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_22),
    .d1(q_12_23),
    .q(q_13_23)
  );
  

  flop_with_mux u_13_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_23),
    .d1(q_12_24),
    .q(q_13_24)
  );
  

  flop_with_mux u_13_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_24),
    .d1(q_12_25),
    .q(q_13_25)
  );
  

  flop_with_mux u_13_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_25),
    .d1(q_12_26),
    .q(q_13_26)
  );
  

  flop_with_mux u_13_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_26),
    .d1(q_12_27),
    .q(q_13_27)
  );
  

  flop_with_mux u_13_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_27),
    .d1(q_12_28),
    .q(q_13_28)
  );
  

  flop_with_mux u_13_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_28),
    .d1(q_12_29),
    .q(q_13_29)
  );
  

  flop_with_mux u_13_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_29),
    .d1(q_12_30),
    .q(q_13_30)
  );
  

  flop_with_mux u_13_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_30),
    .d1(q_12_31),
    .q(q_13_31)
  );
  

  flop_with_mux u_13_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_31),
    .d1(q_12_32),
    .q(q_13_32)
  );
  

  flop_with_mux u_13_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_32),
    .d1(q_12_33),
    .q(q_13_33)
  );
  

  flop_with_mux u_13_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_33),
    .d1(q_12_34),
    .q(q_13_34)
  );
  

  flop_with_mux u_13_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_34),
    .d1(q_12_35),
    .q(q_13_35)
  );
  

  flop_with_mux u_13_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_35),
    .d1(q_12_36),
    .q(q_13_36)
  );
  

  flop_with_mux u_13_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_36),
    .d1(q_12_37),
    .q(q_13_37)
  );
  

  flop_with_mux u_13_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_37),
    .d1(q_12_38),
    .q(q_13_38)
  );
  

  flop_with_mux u_13_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_13_38),
    .d1(q_12_39),
    .q(q_13_39)
  );
  

  flop_with_mux u_14_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_minus1),
    .d1(q_13_0),
    .q(q_14_0)
  );
  

  flop_with_mux u_14_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_0),
    .d1(q_13_1),
    .q(q_14_1)
  );
  

  flop_with_mux u_14_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_1),
    .d1(q_13_2),
    .q(q_14_2)
  );
  

  flop_with_mux u_14_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_2),
    .d1(q_13_3),
    .q(q_14_3)
  );
  

  flop_with_mux u_14_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_3),
    .d1(q_13_4),
    .q(q_14_4)
  );
  

  flop_with_mux u_14_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_4),
    .d1(q_13_5),
    .q(q_14_5)
  );
  

  flop_with_mux u_14_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_5),
    .d1(q_13_6),
    .q(q_14_6)
  );
  

  flop_with_mux u_14_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_6),
    .d1(q_13_7),
    .q(q_14_7)
  );
  

  flop_with_mux u_14_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_7),
    .d1(q_13_8),
    .q(q_14_8)
  );
  

  flop_with_mux u_14_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_8),
    .d1(q_13_9),
    .q(q_14_9)
  );
  

  flop_with_mux u_14_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_9),
    .d1(q_13_10),
    .q(q_14_10)
  );
  

  flop_with_mux u_14_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_10),
    .d1(q_13_11),
    .q(q_14_11)
  );
  

  flop_with_mux u_14_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_11),
    .d1(q_13_12),
    .q(q_14_12)
  );
  

  flop_with_mux u_14_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_12),
    .d1(q_13_13),
    .q(q_14_13)
  );
  

  flop_with_mux u_14_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_13),
    .d1(q_13_14),
    .q(q_14_14)
  );
  

  flop_with_mux u_14_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_14),
    .d1(q_13_15),
    .q(q_14_15)
  );
  

  flop_with_mux u_14_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_15),
    .d1(q_13_16),
    .q(q_14_16)
  );
  

  flop_with_mux u_14_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_16),
    .d1(q_13_17),
    .q(q_14_17)
  );
  

  flop_with_mux u_14_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_17),
    .d1(q_13_18),
    .q(q_14_18)
  );
  

  flop_with_mux u_14_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_18),
    .d1(q_13_19),
    .q(q_14_19)
  );
  

  flop_with_mux u_14_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_19),
    .d1(q_13_20),
    .q(q_14_20)
  );
  

  flop_with_mux u_14_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_20),
    .d1(q_13_21),
    .q(q_14_21)
  );
  

  flop_with_mux u_14_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_21),
    .d1(q_13_22),
    .q(q_14_22)
  );
  

  flop_with_mux u_14_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_22),
    .d1(q_13_23),
    .q(q_14_23)
  );
  

  flop_with_mux u_14_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_23),
    .d1(q_13_24),
    .q(q_14_24)
  );
  

  flop_with_mux u_14_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_24),
    .d1(q_13_25),
    .q(q_14_25)
  );
  

  flop_with_mux u_14_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_25),
    .d1(q_13_26),
    .q(q_14_26)
  );
  

  flop_with_mux u_14_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_26),
    .d1(q_13_27),
    .q(q_14_27)
  );
  

  flop_with_mux u_14_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_27),
    .d1(q_13_28),
    .q(q_14_28)
  );
  

  flop_with_mux u_14_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_28),
    .d1(q_13_29),
    .q(q_14_29)
  );
  

  flop_with_mux u_14_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_29),
    .d1(q_13_30),
    .q(q_14_30)
  );
  

  flop_with_mux u_14_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_30),
    .d1(q_13_31),
    .q(q_14_31)
  );
  

  flop_with_mux u_14_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_31),
    .d1(q_13_32),
    .q(q_14_32)
  );
  

  flop_with_mux u_14_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_32),
    .d1(q_13_33),
    .q(q_14_33)
  );
  

  flop_with_mux u_14_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_33),
    .d1(q_13_34),
    .q(q_14_34)
  );
  

  flop_with_mux u_14_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_34),
    .d1(q_13_35),
    .q(q_14_35)
  );
  

  flop_with_mux u_14_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_35),
    .d1(q_13_36),
    .q(q_14_36)
  );
  

  flop_with_mux u_14_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_36),
    .d1(q_13_37),
    .q(q_14_37)
  );
  

  flop_with_mux u_14_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_37),
    .d1(q_13_38),
    .q(q_14_38)
  );
  

  flop_with_mux u_14_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_14_38),
    .d1(q_13_39),
    .q(q_14_39)
  );
  

  flop_with_mux u_15_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_minus1),
    .d1(q_14_0),
    .q(q_15_0)
  );
  

  flop_with_mux u_15_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_0),
    .d1(q_14_1),
    .q(q_15_1)
  );
  

  flop_with_mux u_15_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_1),
    .d1(q_14_2),
    .q(q_15_2)
  );
  

  flop_with_mux u_15_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_2),
    .d1(q_14_3),
    .q(q_15_3)
  );
  

  flop_with_mux u_15_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_3),
    .d1(q_14_4),
    .q(q_15_4)
  );
  

  flop_with_mux u_15_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_4),
    .d1(q_14_5),
    .q(q_15_5)
  );
  

  flop_with_mux u_15_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_5),
    .d1(q_14_6),
    .q(q_15_6)
  );
  

  flop_with_mux u_15_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_6),
    .d1(q_14_7),
    .q(q_15_7)
  );
  

  flop_with_mux u_15_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_7),
    .d1(q_14_8),
    .q(q_15_8)
  );
  

  flop_with_mux u_15_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_8),
    .d1(q_14_9),
    .q(q_15_9)
  );
  

  flop_with_mux u_15_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_9),
    .d1(q_14_10),
    .q(q_15_10)
  );
  

  flop_with_mux u_15_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_10),
    .d1(q_14_11),
    .q(q_15_11)
  );
  

  flop_with_mux u_15_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_11),
    .d1(q_14_12),
    .q(q_15_12)
  );
  

  flop_with_mux u_15_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_12),
    .d1(q_14_13),
    .q(q_15_13)
  );
  

  flop_with_mux u_15_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_13),
    .d1(q_14_14),
    .q(q_15_14)
  );
  

  flop_with_mux u_15_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_14),
    .d1(q_14_15),
    .q(q_15_15)
  );
  

  flop_with_mux u_15_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_15),
    .d1(q_14_16),
    .q(q_15_16)
  );
  

  flop_with_mux u_15_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_16),
    .d1(q_14_17),
    .q(q_15_17)
  );
  

  flop_with_mux u_15_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_17),
    .d1(q_14_18),
    .q(q_15_18)
  );
  

  flop_with_mux u_15_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_18),
    .d1(q_14_19),
    .q(q_15_19)
  );
  

  flop_with_mux u_15_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_19),
    .d1(q_14_20),
    .q(q_15_20)
  );
  

  flop_with_mux u_15_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_20),
    .d1(q_14_21),
    .q(q_15_21)
  );
  

  flop_with_mux u_15_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_21),
    .d1(q_14_22),
    .q(q_15_22)
  );
  

  flop_with_mux u_15_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_22),
    .d1(q_14_23),
    .q(q_15_23)
  );
  

  flop_with_mux u_15_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_23),
    .d1(q_14_24),
    .q(q_15_24)
  );
  

  flop_with_mux u_15_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_24),
    .d1(q_14_25),
    .q(q_15_25)
  );
  

  flop_with_mux u_15_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_25),
    .d1(q_14_26),
    .q(q_15_26)
  );
  

  flop_with_mux u_15_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_26),
    .d1(q_14_27),
    .q(q_15_27)
  );
  

  flop_with_mux u_15_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_27),
    .d1(q_14_28),
    .q(q_15_28)
  );
  

  flop_with_mux u_15_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_28),
    .d1(q_14_29),
    .q(q_15_29)
  );
  

  flop_with_mux u_15_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_29),
    .d1(q_14_30),
    .q(q_15_30)
  );
  

  flop_with_mux u_15_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_30),
    .d1(q_14_31),
    .q(q_15_31)
  );
  

  flop_with_mux u_15_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_31),
    .d1(q_14_32),
    .q(q_15_32)
  );
  

  flop_with_mux u_15_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_32),
    .d1(q_14_33),
    .q(q_15_33)
  );
  

  flop_with_mux u_15_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_33),
    .d1(q_14_34),
    .q(q_15_34)
  );
  

  flop_with_mux u_15_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_34),
    .d1(q_14_35),
    .q(q_15_35)
  );
  

  flop_with_mux u_15_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_35),
    .d1(q_14_36),
    .q(q_15_36)
  );
  

  flop_with_mux u_15_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_36),
    .d1(q_14_37),
    .q(q_15_37)
  );
  

  flop_with_mux u_15_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_37),
    .d1(q_14_38),
    .q(q_15_38)
  );
  

  flop_with_mux u_15_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_15_38),
    .d1(q_14_39),
    .q(q_15_39)
  );
  

  flop_with_mux u_16_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_minus1),
    .d1(q_15_0),
    .q(q_16_0)
  );
  

  flop_with_mux u_16_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_0),
    .d1(q_15_1),
    .q(q_16_1)
  );
  

  flop_with_mux u_16_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_1),
    .d1(q_15_2),
    .q(q_16_2)
  );
  

  flop_with_mux u_16_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_2),
    .d1(q_15_3),
    .q(q_16_3)
  );
  

  flop_with_mux u_16_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_3),
    .d1(q_15_4),
    .q(q_16_4)
  );
  

  flop_with_mux u_16_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_4),
    .d1(q_15_5),
    .q(q_16_5)
  );
  

  flop_with_mux u_16_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_5),
    .d1(q_15_6),
    .q(q_16_6)
  );
  

  flop_with_mux u_16_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_6),
    .d1(q_15_7),
    .q(q_16_7)
  );
  

  flop_with_mux u_16_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_7),
    .d1(q_15_8),
    .q(q_16_8)
  );
  

  flop_with_mux u_16_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_8),
    .d1(q_15_9),
    .q(q_16_9)
  );
  

  flop_with_mux u_16_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_9),
    .d1(q_15_10),
    .q(q_16_10)
  );
  

  flop_with_mux u_16_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_10),
    .d1(q_15_11),
    .q(q_16_11)
  );
  

  flop_with_mux u_16_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_11),
    .d1(q_15_12),
    .q(q_16_12)
  );
  

  flop_with_mux u_16_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_12),
    .d1(q_15_13),
    .q(q_16_13)
  );
  

  flop_with_mux u_16_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_13),
    .d1(q_15_14),
    .q(q_16_14)
  );
  

  flop_with_mux u_16_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_14),
    .d1(q_15_15),
    .q(q_16_15)
  );
  

  flop_with_mux u_16_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_15),
    .d1(q_15_16),
    .q(q_16_16)
  );
  

  flop_with_mux u_16_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_16),
    .d1(q_15_17),
    .q(q_16_17)
  );
  

  flop_with_mux u_16_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_17),
    .d1(q_15_18),
    .q(q_16_18)
  );
  

  flop_with_mux u_16_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_18),
    .d1(q_15_19),
    .q(q_16_19)
  );
  

  flop_with_mux u_16_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_19),
    .d1(q_15_20),
    .q(q_16_20)
  );
  

  flop_with_mux u_16_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_20),
    .d1(q_15_21),
    .q(q_16_21)
  );
  

  flop_with_mux u_16_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_21),
    .d1(q_15_22),
    .q(q_16_22)
  );
  

  flop_with_mux u_16_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_22),
    .d1(q_15_23),
    .q(q_16_23)
  );
  

  flop_with_mux u_16_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_23),
    .d1(q_15_24),
    .q(q_16_24)
  );
  

  flop_with_mux u_16_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_24),
    .d1(q_15_25),
    .q(q_16_25)
  );
  

  flop_with_mux u_16_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_25),
    .d1(q_15_26),
    .q(q_16_26)
  );
  

  flop_with_mux u_16_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_26),
    .d1(q_15_27),
    .q(q_16_27)
  );
  

  flop_with_mux u_16_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_27),
    .d1(q_15_28),
    .q(q_16_28)
  );
  

  flop_with_mux u_16_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_28),
    .d1(q_15_29),
    .q(q_16_29)
  );
  

  flop_with_mux u_16_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_29),
    .d1(q_15_30),
    .q(q_16_30)
  );
  

  flop_with_mux u_16_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_30),
    .d1(q_15_31),
    .q(q_16_31)
  );
  

  flop_with_mux u_16_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_31),
    .d1(q_15_32),
    .q(q_16_32)
  );
  

  flop_with_mux u_16_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_32),
    .d1(q_15_33),
    .q(q_16_33)
  );
  

  flop_with_mux u_16_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_33),
    .d1(q_15_34),
    .q(q_16_34)
  );
  

  flop_with_mux u_16_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_34),
    .d1(q_15_35),
    .q(q_16_35)
  );
  

  flop_with_mux u_16_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_35),
    .d1(q_15_36),
    .q(q_16_36)
  );
  

  flop_with_mux u_16_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_36),
    .d1(q_15_37),
    .q(q_16_37)
  );
  

  flop_with_mux u_16_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_37),
    .d1(q_15_38),
    .q(q_16_38)
  );
  

  flop_with_mux u_16_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_16_38),
    .d1(q_15_39),
    .q(q_16_39)
  );
  

  flop_with_mux u_17_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_minus1),
    .d1(q_16_0),
    .q(q_17_0)
  );
  

  flop_with_mux u_17_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_0),
    .d1(q_16_1),
    .q(q_17_1)
  );
  

  flop_with_mux u_17_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_1),
    .d1(q_16_2),
    .q(q_17_2)
  );
  

  flop_with_mux u_17_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_2),
    .d1(q_16_3),
    .q(q_17_3)
  );
  

  flop_with_mux u_17_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_3),
    .d1(q_16_4),
    .q(q_17_4)
  );
  

  flop_with_mux u_17_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_4),
    .d1(q_16_5),
    .q(q_17_5)
  );
  

  flop_with_mux u_17_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_5),
    .d1(q_16_6),
    .q(q_17_6)
  );
  

  flop_with_mux u_17_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_6),
    .d1(q_16_7),
    .q(q_17_7)
  );
  

  flop_with_mux u_17_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_7),
    .d1(q_16_8),
    .q(q_17_8)
  );
  

  flop_with_mux u_17_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_8),
    .d1(q_16_9),
    .q(q_17_9)
  );
  

  flop_with_mux u_17_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_9),
    .d1(q_16_10),
    .q(q_17_10)
  );
  

  flop_with_mux u_17_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_10),
    .d1(q_16_11),
    .q(q_17_11)
  );
  

  flop_with_mux u_17_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_11),
    .d1(q_16_12),
    .q(q_17_12)
  );
  

  flop_with_mux u_17_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_12),
    .d1(q_16_13),
    .q(q_17_13)
  );
  

  flop_with_mux u_17_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_13),
    .d1(q_16_14),
    .q(q_17_14)
  );
  

  flop_with_mux u_17_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_14),
    .d1(q_16_15),
    .q(q_17_15)
  );
  

  flop_with_mux u_17_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_15),
    .d1(q_16_16),
    .q(q_17_16)
  );
  

  flop_with_mux u_17_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_16),
    .d1(q_16_17),
    .q(q_17_17)
  );
  

  flop_with_mux u_17_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_17),
    .d1(q_16_18),
    .q(q_17_18)
  );
  

  flop_with_mux u_17_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_18),
    .d1(q_16_19),
    .q(q_17_19)
  );
  

  flop_with_mux u_17_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_19),
    .d1(q_16_20),
    .q(q_17_20)
  );
  

  flop_with_mux u_17_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_20),
    .d1(q_16_21),
    .q(q_17_21)
  );
  

  flop_with_mux u_17_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_21),
    .d1(q_16_22),
    .q(q_17_22)
  );
  

  flop_with_mux u_17_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_22),
    .d1(q_16_23),
    .q(q_17_23)
  );
  

  flop_with_mux u_17_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_23),
    .d1(q_16_24),
    .q(q_17_24)
  );
  

  flop_with_mux u_17_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_24),
    .d1(q_16_25),
    .q(q_17_25)
  );
  

  flop_with_mux u_17_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_25),
    .d1(q_16_26),
    .q(q_17_26)
  );
  

  flop_with_mux u_17_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_26),
    .d1(q_16_27),
    .q(q_17_27)
  );
  

  flop_with_mux u_17_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_27),
    .d1(q_16_28),
    .q(q_17_28)
  );
  

  flop_with_mux u_17_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_28),
    .d1(q_16_29),
    .q(q_17_29)
  );
  

  flop_with_mux u_17_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_29),
    .d1(q_16_30),
    .q(q_17_30)
  );
  

  flop_with_mux u_17_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_30),
    .d1(q_16_31),
    .q(q_17_31)
  );
  

  flop_with_mux u_17_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_31),
    .d1(q_16_32),
    .q(q_17_32)
  );
  

  flop_with_mux u_17_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_32),
    .d1(q_16_33),
    .q(q_17_33)
  );
  

  flop_with_mux u_17_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_33),
    .d1(q_16_34),
    .q(q_17_34)
  );
  

  flop_with_mux u_17_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_34),
    .d1(q_16_35),
    .q(q_17_35)
  );
  

  flop_with_mux u_17_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_35),
    .d1(q_16_36),
    .q(q_17_36)
  );
  

  flop_with_mux u_17_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_36),
    .d1(q_16_37),
    .q(q_17_37)
  );
  

  flop_with_mux u_17_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_37),
    .d1(q_16_38),
    .q(q_17_38)
  );
  

  flop_with_mux u_17_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_17_38),
    .d1(q_16_39),
    .q(q_17_39)
  );
  

  flop_with_mux u_18_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_minus1),
    .d1(q_17_0),
    .q(q_18_0)
  );
  

  flop_with_mux u_18_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_0),
    .d1(q_17_1),
    .q(q_18_1)
  );
  

  flop_with_mux u_18_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_1),
    .d1(q_17_2),
    .q(q_18_2)
  );
  

  flop_with_mux u_18_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_2),
    .d1(q_17_3),
    .q(q_18_3)
  );
  

  flop_with_mux u_18_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_3),
    .d1(q_17_4),
    .q(q_18_4)
  );
  

  flop_with_mux u_18_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_4),
    .d1(q_17_5),
    .q(q_18_5)
  );
  

  flop_with_mux u_18_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_5),
    .d1(q_17_6),
    .q(q_18_6)
  );
  

  flop_with_mux u_18_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_6),
    .d1(q_17_7),
    .q(q_18_7)
  );
  

  flop_with_mux u_18_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_7),
    .d1(q_17_8),
    .q(q_18_8)
  );
  

  flop_with_mux u_18_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_8),
    .d1(q_17_9),
    .q(q_18_9)
  );
  

  flop_with_mux u_18_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_9),
    .d1(q_17_10),
    .q(q_18_10)
  );
  

  flop_with_mux u_18_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_10),
    .d1(q_17_11),
    .q(q_18_11)
  );
  

  flop_with_mux u_18_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_11),
    .d1(q_17_12),
    .q(q_18_12)
  );
  

  flop_with_mux u_18_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_12),
    .d1(q_17_13),
    .q(q_18_13)
  );
  

  flop_with_mux u_18_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_13),
    .d1(q_17_14),
    .q(q_18_14)
  );
  

  flop_with_mux u_18_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_14),
    .d1(q_17_15),
    .q(q_18_15)
  );
  

  flop_with_mux u_18_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_15),
    .d1(q_17_16),
    .q(q_18_16)
  );
  

  flop_with_mux u_18_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_16),
    .d1(q_17_17),
    .q(q_18_17)
  );
  

  flop_with_mux u_18_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_17),
    .d1(q_17_18),
    .q(q_18_18)
  );
  

  flop_with_mux u_18_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_18),
    .d1(q_17_19),
    .q(q_18_19)
  );
  

  flop_with_mux u_18_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_19),
    .d1(q_17_20),
    .q(q_18_20)
  );
  

  flop_with_mux u_18_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_20),
    .d1(q_17_21),
    .q(q_18_21)
  );
  

  flop_with_mux u_18_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_21),
    .d1(q_17_22),
    .q(q_18_22)
  );
  

  flop_with_mux u_18_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_22),
    .d1(q_17_23),
    .q(q_18_23)
  );
  

  flop_with_mux u_18_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_23),
    .d1(q_17_24),
    .q(q_18_24)
  );
  

  flop_with_mux u_18_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_24),
    .d1(q_17_25),
    .q(q_18_25)
  );
  

  flop_with_mux u_18_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_25),
    .d1(q_17_26),
    .q(q_18_26)
  );
  

  flop_with_mux u_18_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_26),
    .d1(q_17_27),
    .q(q_18_27)
  );
  

  flop_with_mux u_18_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_27),
    .d1(q_17_28),
    .q(q_18_28)
  );
  

  flop_with_mux u_18_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_28),
    .d1(q_17_29),
    .q(q_18_29)
  );
  

  flop_with_mux u_18_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_29),
    .d1(q_17_30),
    .q(q_18_30)
  );
  

  flop_with_mux u_18_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_30),
    .d1(q_17_31),
    .q(q_18_31)
  );
  

  flop_with_mux u_18_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_31),
    .d1(q_17_32),
    .q(q_18_32)
  );
  

  flop_with_mux u_18_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_32),
    .d1(q_17_33),
    .q(q_18_33)
  );
  

  flop_with_mux u_18_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_33),
    .d1(q_17_34),
    .q(q_18_34)
  );
  

  flop_with_mux u_18_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_34),
    .d1(q_17_35),
    .q(q_18_35)
  );
  

  flop_with_mux u_18_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_35),
    .d1(q_17_36),
    .q(q_18_36)
  );
  

  flop_with_mux u_18_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_36),
    .d1(q_17_37),
    .q(q_18_37)
  );
  

  flop_with_mux u_18_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_37),
    .d1(q_17_38),
    .q(q_18_38)
  );
  

  flop_with_mux u_18_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_18_38),
    .d1(q_17_39),
    .q(q_18_39)
  );
  

  flop_with_mux u_19_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_minus1),
    .d1(q_18_0),
    .q(q_19_0)
  );
  

  flop_with_mux u_19_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_0),
    .d1(q_18_1),
    .q(q_19_1)
  );
  

  flop_with_mux u_19_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_1),
    .d1(q_18_2),
    .q(q_19_2)
  );
  

  flop_with_mux u_19_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_2),
    .d1(q_18_3),
    .q(q_19_3)
  );
  

  flop_with_mux u_19_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_3),
    .d1(q_18_4),
    .q(q_19_4)
  );
  

  flop_with_mux u_19_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_4),
    .d1(q_18_5),
    .q(q_19_5)
  );
  

  flop_with_mux u_19_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_5),
    .d1(q_18_6),
    .q(q_19_6)
  );
  

  flop_with_mux u_19_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_6),
    .d1(q_18_7),
    .q(q_19_7)
  );
  

  flop_with_mux u_19_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_7),
    .d1(q_18_8),
    .q(q_19_8)
  );
  

  flop_with_mux u_19_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_8),
    .d1(q_18_9),
    .q(q_19_9)
  );
  

  flop_with_mux u_19_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_9),
    .d1(q_18_10),
    .q(q_19_10)
  );
  

  flop_with_mux u_19_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_10),
    .d1(q_18_11),
    .q(q_19_11)
  );
  

  flop_with_mux u_19_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_11),
    .d1(q_18_12),
    .q(q_19_12)
  );
  

  flop_with_mux u_19_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_12),
    .d1(q_18_13),
    .q(q_19_13)
  );
  

  flop_with_mux u_19_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_13),
    .d1(q_18_14),
    .q(q_19_14)
  );
  

  flop_with_mux u_19_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_14),
    .d1(q_18_15),
    .q(q_19_15)
  );
  

  flop_with_mux u_19_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_15),
    .d1(q_18_16),
    .q(q_19_16)
  );
  

  flop_with_mux u_19_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_16),
    .d1(q_18_17),
    .q(q_19_17)
  );
  

  flop_with_mux u_19_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_17),
    .d1(q_18_18),
    .q(q_19_18)
  );
  

  flop_with_mux u_19_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_18),
    .d1(q_18_19),
    .q(q_19_19)
  );
  

  flop_with_mux u_19_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_19),
    .d1(q_18_20),
    .q(q_19_20)
  );
  

  flop_with_mux u_19_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_20),
    .d1(q_18_21),
    .q(q_19_21)
  );
  

  flop_with_mux u_19_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_21),
    .d1(q_18_22),
    .q(q_19_22)
  );
  

  flop_with_mux u_19_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_22),
    .d1(q_18_23),
    .q(q_19_23)
  );
  

  flop_with_mux u_19_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_23),
    .d1(q_18_24),
    .q(q_19_24)
  );
  

  flop_with_mux u_19_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_24),
    .d1(q_18_25),
    .q(q_19_25)
  );
  

  flop_with_mux u_19_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_25),
    .d1(q_18_26),
    .q(q_19_26)
  );
  

  flop_with_mux u_19_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_26),
    .d1(q_18_27),
    .q(q_19_27)
  );
  

  flop_with_mux u_19_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_27),
    .d1(q_18_28),
    .q(q_19_28)
  );
  

  flop_with_mux u_19_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_28),
    .d1(q_18_29),
    .q(q_19_29)
  );
  

  flop_with_mux u_19_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_29),
    .d1(q_18_30),
    .q(q_19_30)
  );
  

  flop_with_mux u_19_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_30),
    .d1(q_18_31),
    .q(q_19_31)
  );
  

  flop_with_mux u_19_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_31),
    .d1(q_18_32),
    .q(q_19_32)
  );
  

  flop_with_mux u_19_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_32),
    .d1(q_18_33),
    .q(q_19_33)
  );
  

  flop_with_mux u_19_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_33),
    .d1(q_18_34),
    .q(q_19_34)
  );
  

  flop_with_mux u_19_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_34),
    .d1(q_18_35),
    .q(q_19_35)
  );
  

  flop_with_mux u_19_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_35),
    .d1(q_18_36),
    .q(q_19_36)
  );
  

  flop_with_mux u_19_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_36),
    .d1(q_18_37),
    .q(q_19_37)
  );
  

  flop_with_mux u_19_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_37),
    .d1(q_18_38),
    .q(q_19_38)
  );
  

  flop_with_mux u_19_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_19_38),
    .d1(q_18_39),
    .q(q_19_39)
  );
  

  flop_with_mux u_20_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_minus1),
    .d1(q_19_0),
    .q(q_20_0)
  );
  

  flop_with_mux u_20_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_0),
    .d1(q_19_1),
    .q(q_20_1)
  );
  

  flop_with_mux u_20_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_1),
    .d1(q_19_2),
    .q(q_20_2)
  );
  

  flop_with_mux u_20_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_2),
    .d1(q_19_3),
    .q(q_20_3)
  );
  

  flop_with_mux u_20_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_3),
    .d1(q_19_4),
    .q(q_20_4)
  );
  

  flop_with_mux u_20_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_4),
    .d1(q_19_5),
    .q(q_20_5)
  );
  

  flop_with_mux u_20_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_5),
    .d1(q_19_6),
    .q(q_20_6)
  );
  

  flop_with_mux u_20_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_6),
    .d1(q_19_7),
    .q(q_20_7)
  );
  

  flop_with_mux u_20_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_7),
    .d1(q_19_8),
    .q(q_20_8)
  );
  

  flop_with_mux u_20_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_8),
    .d1(q_19_9),
    .q(q_20_9)
  );
  

  flop_with_mux u_20_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_9),
    .d1(q_19_10),
    .q(q_20_10)
  );
  

  flop_with_mux u_20_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_10),
    .d1(q_19_11),
    .q(q_20_11)
  );
  

  flop_with_mux u_20_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_11),
    .d1(q_19_12),
    .q(q_20_12)
  );
  

  flop_with_mux u_20_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_12),
    .d1(q_19_13),
    .q(q_20_13)
  );
  

  flop_with_mux u_20_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_13),
    .d1(q_19_14),
    .q(q_20_14)
  );
  

  flop_with_mux u_20_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_14),
    .d1(q_19_15),
    .q(q_20_15)
  );
  

  flop_with_mux u_20_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_15),
    .d1(q_19_16),
    .q(q_20_16)
  );
  

  flop_with_mux u_20_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_16),
    .d1(q_19_17),
    .q(q_20_17)
  );
  

  flop_with_mux u_20_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_17),
    .d1(q_19_18),
    .q(q_20_18)
  );
  

  flop_with_mux u_20_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_18),
    .d1(q_19_19),
    .q(q_20_19)
  );
  

  flop_with_mux u_20_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_19),
    .d1(q_19_20),
    .q(q_20_20)
  );
  

  flop_with_mux u_20_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_20),
    .d1(q_19_21),
    .q(q_20_21)
  );
  

  flop_with_mux u_20_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_21),
    .d1(q_19_22),
    .q(q_20_22)
  );
  

  flop_with_mux u_20_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_22),
    .d1(q_19_23),
    .q(q_20_23)
  );
  

  flop_with_mux u_20_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_23),
    .d1(q_19_24),
    .q(q_20_24)
  );
  

  flop_with_mux u_20_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_24),
    .d1(q_19_25),
    .q(q_20_25)
  );
  

  flop_with_mux u_20_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_25),
    .d1(q_19_26),
    .q(q_20_26)
  );
  

  flop_with_mux u_20_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_26),
    .d1(q_19_27),
    .q(q_20_27)
  );
  

  flop_with_mux u_20_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_27),
    .d1(q_19_28),
    .q(q_20_28)
  );
  

  flop_with_mux u_20_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_28),
    .d1(q_19_29),
    .q(q_20_29)
  );
  

  flop_with_mux u_20_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_29),
    .d1(q_19_30),
    .q(q_20_30)
  );
  

  flop_with_mux u_20_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_30),
    .d1(q_19_31),
    .q(q_20_31)
  );
  

  flop_with_mux u_20_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_31),
    .d1(q_19_32),
    .q(q_20_32)
  );
  

  flop_with_mux u_20_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_32),
    .d1(q_19_33),
    .q(q_20_33)
  );
  

  flop_with_mux u_20_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_33),
    .d1(q_19_34),
    .q(q_20_34)
  );
  

  flop_with_mux u_20_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_34),
    .d1(q_19_35),
    .q(q_20_35)
  );
  

  flop_with_mux u_20_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_35),
    .d1(q_19_36),
    .q(q_20_36)
  );
  

  flop_with_mux u_20_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_36),
    .d1(q_19_37),
    .q(q_20_37)
  );
  

  flop_with_mux u_20_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_37),
    .d1(q_19_38),
    .q(q_20_38)
  );
  

  flop_with_mux u_20_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_20_38),
    .d1(q_19_39),
    .q(q_20_39)
  );
  

  flop_with_mux u_21_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_minus1),
    .d1(q_20_0),
    .q(q_21_0)
  );
  

  flop_with_mux u_21_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_0),
    .d1(q_20_1),
    .q(q_21_1)
  );
  

  flop_with_mux u_21_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_1),
    .d1(q_20_2),
    .q(q_21_2)
  );
  

  flop_with_mux u_21_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_2),
    .d1(q_20_3),
    .q(q_21_3)
  );
  

  flop_with_mux u_21_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_3),
    .d1(q_20_4),
    .q(q_21_4)
  );
  

  flop_with_mux u_21_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_4),
    .d1(q_20_5),
    .q(q_21_5)
  );
  

  flop_with_mux u_21_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_5),
    .d1(q_20_6),
    .q(q_21_6)
  );
  

  flop_with_mux u_21_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_6),
    .d1(q_20_7),
    .q(q_21_7)
  );
  

  flop_with_mux u_21_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_7),
    .d1(q_20_8),
    .q(q_21_8)
  );
  

  flop_with_mux u_21_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_8),
    .d1(q_20_9),
    .q(q_21_9)
  );
  

  flop_with_mux u_21_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_9),
    .d1(q_20_10),
    .q(q_21_10)
  );
  

  flop_with_mux u_21_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_10),
    .d1(q_20_11),
    .q(q_21_11)
  );
  

  flop_with_mux u_21_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_11),
    .d1(q_20_12),
    .q(q_21_12)
  );
  

  flop_with_mux u_21_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_12),
    .d1(q_20_13),
    .q(q_21_13)
  );
  

  flop_with_mux u_21_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_13),
    .d1(q_20_14),
    .q(q_21_14)
  );
  

  flop_with_mux u_21_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_14),
    .d1(q_20_15),
    .q(q_21_15)
  );
  

  flop_with_mux u_21_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_15),
    .d1(q_20_16),
    .q(q_21_16)
  );
  

  flop_with_mux u_21_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_16),
    .d1(q_20_17),
    .q(q_21_17)
  );
  

  flop_with_mux u_21_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_17),
    .d1(q_20_18),
    .q(q_21_18)
  );
  

  flop_with_mux u_21_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_18),
    .d1(q_20_19),
    .q(q_21_19)
  );
  

  flop_with_mux u_21_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_19),
    .d1(q_20_20),
    .q(q_21_20)
  );
  

  flop_with_mux u_21_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_20),
    .d1(q_20_21),
    .q(q_21_21)
  );
  

  flop_with_mux u_21_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_21),
    .d1(q_20_22),
    .q(q_21_22)
  );
  

  flop_with_mux u_21_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_22),
    .d1(q_20_23),
    .q(q_21_23)
  );
  

  flop_with_mux u_21_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_23),
    .d1(q_20_24),
    .q(q_21_24)
  );
  

  flop_with_mux u_21_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_24),
    .d1(q_20_25),
    .q(q_21_25)
  );
  

  flop_with_mux u_21_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_25),
    .d1(q_20_26),
    .q(q_21_26)
  );
  

  flop_with_mux u_21_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_26),
    .d1(q_20_27),
    .q(q_21_27)
  );
  

  flop_with_mux u_21_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_27),
    .d1(q_20_28),
    .q(q_21_28)
  );
  

  flop_with_mux u_21_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_28),
    .d1(q_20_29),
    .q(q_21_29)
  );
  

  flop_with_mux u_21_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_29),
    .d1(q_20_30),
    .q(q_21_30)
  );
  

  flop_with_mux u_21_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_30),
    .d1(q_20_31),
    .q(q_21_31)
  );
  

  flop_with_mux u_21_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_31),
    .d1(q_20_32),
    .q(q_21_32)
  );
  

  flop_with_mux u_21_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_32),
    .d1(q_20_33),
    .q(q_21_33)
  );
  

  flop_with_mux u_21_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_33),
    .d1(q_20_34),
    .q(q_21_34)
  );
  

  flop_with_mux u_21_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_34),
    .d1(q_20_35),
    .q(q_21_35)
  );
  

  flop_with_mux u_21_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_35),
    .d1(q_20_36),
    .q(q_21_36)
  );
  

  flop_with_mux u_21_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_36),
    .d1(q_20_37),
    .q(q_21_37)
  );
  

  flop_with_mux u_21_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_37),
    .d1(q_20_38),
    .q(q_21_38)
  );
  

  flop_with_mux u_21_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_21_38),
    .d1(q_20_39),
    .q(q_21_39)
  );
  

  flop_with_mux u_22_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_minus1),
    .d1(q_21_0),
    .q(q_22_0)
  );
  

  flop_with_mux u_22_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_0),
    .d1(q_21_1),
    .q(q_22_1)
  );
  

  flop_with_mux u_22_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_1),
    .d1(q_21_2),
    .q(q_22_2)
  );
  

  flop_with_mux u_22_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_2),
    .d1(q_21_3),
    .q(q_22_3)
  );
  

  flop_with_mux u_22_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_3),
    .d1(q_21_4),
    .q(q_22_4)
  );
  

  flop_with_mux u_22_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_4),
    .d1(q_21_5),
    .q(q_22_5)
  );
  

  flop_with_mux u_22_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_5),
    .d1(q_21_6),
    .q(q_22_6)
  );
  

  flop_with_mux u_22_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_6),
    .d1(q_21_7),
    .q(q_22_7)
  );
  

  flop_with_mux u_22_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_7),
    .d1(q_21_8),
    .q(q_22_8)
  );
  

  flop_with_mux u_22_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_8),
    .d1(q_21_9),
    .q(q_22_9)
  );
  

  flop_with_mux u_22_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_9),
    .d1(q_21_10),
    .q(q_22_10)
  );
  

  flop_with_mux u_22_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_10),
    .d1(q_21_11),
    .q(q_22_11)
  );
  

  flop_with_mux u_22_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_11),
    .d1(q_21_12),
    .q(q_22_12)
  );
  

  flop_with_mux u_22_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_12),
    .d1(q_21_13),
    .q(q_22_13)
  );
  

  flop_with_mux u_22_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_13),
    .d1(q_21_14),
    .q(q_22_14)
  );
  

  flop_with_mux u_22_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_14),
    .d1(q_21_15),
    .q(q_22_15)
  );
  

  flop_with_mux u_22_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_15),
    .d1(q_21_16),
    .q(q_22_16)
  );
  

  flop_with_mux u_22_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_16),
    .d1(q_21_17),
    .q(q_22_17)
  );
  

  flop_with_mux u_22_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_17),
    .d1(q_21_18),
    .q(q_22_18)
  );
  

  flop_with_mux u_22_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_18),
    .d1(q_21_19),
    .q(q_22_19)
  );
  

  flop_with_mux u_22_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_19),
    .d1(q_21_20),
    .q(q_22_20)
  );
  

  flop_with_mux u_22_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_20),
    .d1(q_21_21),
    .q(q_22_21)
  );
  

  flop_with_mux u_22_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_21),
    .d1(q_21_22),
    .q(q_22_22)
  );
  

  flop_with_mux u_22_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_22),
    .d1(q_21_23),
    .q(q_22_23)
  );
  

  flop_with_mux u_22_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_23),
    .d1(q_21_24),
    .q(q_22_24)
  );
  

  flop_with_mux u_22_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_24),
    .d1(q_21_25),
    .q(q_22_25)
  );
  

  flop_with_mux u_22_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_25),
    .d1(q_21_26),
    .q(q_22_26)
  );
  

  flop_with_mux u_22_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_26),
    .d1(q_21_27),
    .q(q_22_27)
  );
  

  flop_with_mux u_22_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_27),
    .d1(q_21_28),
    .q(q_22_28)
  );
  

  flop_with_mux u_22_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_28),
    .d1(q_21_29),
    .q(q_22_29)
  );
  

  flop_with_mux u_22_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_29),
    .d1(q_21_30),
    .q(q_22_30)
  );
  

  flop_with_mux u_22_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_30),
    .d1(q_21_31),
    .q(q_22_31)
  );
  

  flop_with_mux u_22_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_31),
    .d1(q_21_32),
    .q(q_22_32)
  );
  

  flop_with_mux u_22_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_32),
    .d1(q_21_33),
    .q(q_22_33)
  );
  

  flop_with_mux u_22_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_33),
    .d1(q_21_34),
    .q(q_22_34)
  );
  

  flop_with_mux u_22_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_34),
    .d1(q_21_35),
    .q(q_22_35)
  );
  

  flop_with_mux u_22_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_35),
    .d1(q_21_36),
    .q(q_22_36)
  );
  

  flop_with_mux u_22_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_36),
    .d1(q_21_37),
    .q(q_22_37)
  );
  

  flop_with_mux u_22_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_37),
    .d1(q_21_38),
    .q(q_22_38)
  );
  

  flop_with_mux u_22_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_22_38),
    .d1(q_21_39),
    .q(q_22_39)
  );
  

  flop_with_mux u_23_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_minus1),
    .d1(q_22_0),
    .q(q_23_0)
  );
  

  flop_with_mux u_23_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_0),
    .d1(q_22_1),
    .q(q_23_1)
  );
  

  flop_with_mux u_23_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_1),
    .d1(q_22_2),
    .q(q_23_2)
  );
  

  flop_with_mux u_23_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_2),
    .d1(q_22_3),
    .q(q_23_3)
  );
  

  flop_with_mux u_23_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_3),
    .d1(q_22_4),
    .q(q_23_4)
  );
  

  flop_with_mux u_23_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_4),
    .d1(q_22_5),
    .q(q_23_5)
  );
  

  flop_with_mux u_23_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_5),
    .d1(q_22_6),
    .q(q_23_6)
  );
  

  flop_with_mux u_23_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_6),
    .d1(q_22_7),
    .q(q_23_7)
  );
  

  flop_with_mux u_23_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_7),
    .d1(q_22_8),
    .q(q_23_8)
  );
  

  flop_with_mux u_23_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_8),
    .d1(q_22_9),
    .q(q_23_9)
  );
  

  flop_with_mux u_23_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_9),
    .d1(q_22_10),
    .q(q_23_10)
  );
  

  flop_with_mux u_23_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_10),
    .d1(q_22_11),
    .q(q_23_11)
  );
  

  flop_with_mux u_23_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_11),
    .d1(q_22_12),
    .q(q_23_12)
  );
  

  flop_with_mux u_23_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_12),
    .d1(q_22_13),
    .q(q_23_13)
  );
  

  flop_with_mux u_23_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_13),
    .d1(q_22_14),
    .q(q_23_14)
  );
  

  flop_with_mux u_23_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_14),
    .d1(q_22_15),
    .q(q_23_15)
  );
  

  flop_with_mux u_23_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_15),
    .d1(q_22_16),
    .q(q_23_16)
  );
  

  flop_with_mux u_23_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_16),
    .d1(q_22_17),
    .q(q_23_17)
  );
  

  flop_with_mux u_23_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_17),
    .d1(q_22_18),
    .q(q_23_18)
  );
  

  flop_with_mux u_23_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_18),
    .d1(q_22_19),
    .q(q_23_19)
  );
  

  flop_with_mux u_23_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_19),
    .d1(q_22_20),
    .q(q_23_20)
  );
  

  flop_with_mux u_23_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_20),
    .d1(q_22_21),
    .q(q_23_21)
  );
  

  flop_with_mux u_23_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_21),
    .d1(q_22_22),
    .q(q_23_22)
  );
  

  flop_with_mux u_23_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_22),
    .d1(q_22_23),
    .q(q_23_23)
  );
  

  flop_with_mux u_23_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_23),
    .d1(q_22_24),
    .q(q_23_24)
  );
  

  flop_with_mux u_23_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_24),
    .d1(q_22_25),
    .q(q_23_25)
  );
  

  flop_with_mux u_23_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_25),
    .d1(q_22_26),
    .q(q_23_26)
  );
  

  flop_with_mux u_23_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_26),
    .d1(q_22_27),
    .q(q_23_27)
  );
  

  flop_with_mux u_23_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_27),
    .d1(q_22_28),
    .q(q_23_28)
  );
  

  flop_with_mux u_23_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_28),
    .d1(q_22_29),
    .q(q_23_29)
  );
  

  flop_with_mux u_23_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_29),
    .d1(q_22_30),
    .q(q_23_30)
  );
  

  flop_with_mux u_23_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_30),
    .d1(q_22_31),
    .q(q_23_31)
  );
  

  flop_with_mux u_23_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_31),
    .d1(q_22_32),
    .q(q_23_32)
  );
  

  flop_with_mux u_23_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_32),
    .d1(q_22_33),
    .q(q_23_33)
  );
  

  flop_with_mux u_23_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_33),
    .d1(q_22_34),
    .q(q_23_34)
  );
  

  flop_with_mux u_23_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_34),
    .d1(q_22_35),
    .q(q_23_35)
  );
  

  flop_with_mux u_23_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_35),
    .d1(q_22_36),
    .q(q_23_36)
  );
  

  flop_with_mux u_23_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_36),
    .d1(q_22_37),
    .q(q_23_37)
  );
  

  flop_with_mux u_23_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_37),
    .d1(q_22_38),
    .q(q_23_38)
  );
  

  flop_with_mux u_23_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_23_38),
    .d1(q_22_39),
    .q(q_23_39)
  );
  

  flop_with_mux u_24_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_minus1),
    .d1(q_23_0),
    .q(q_24_0)
  );
  

  flop_with_mux u_24_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_0),
    .d1(q_23_1),
    .q(q_24_1)
  );
  

  flop_with_mux u_24_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_1),
    .d1(q_23_2),
    .q(q_24_2)
  );
  

  flop_with_mux u_24_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_2),
    .d1(q_23_3),
    .q(q_24_3)
  );
  

  flop_with_mux u_24_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_3),
    .d1(q_23_4),
    .q(q_24_4)
  );
  

  flop_with_mux u_24_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_4),
    .d1(q_23_5),
    .q(q_24_5)
  );
  

  flop_with_mux u_24_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_5),
    .d1(q_23_6),
    .q(q_24_6)
  );
  

  flop_with_mux u_24_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_6),
    .d1(q_23_7),
    .q(q_24_7)
  );
  

  flop_with_mux u_24_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_7),
    .d1(q_23_8),
    .q(q_24_8)
  );
  

  flop_with_mux u_24_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_8),
    .d1(q_23_9),
    .q(q_24_9)
  );
  

  flop_with_mux u_24_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_9),
    .d1(q_23_10),
    .q(q_24_10)
  );
  

  flop_with_mux u_24_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_10),
    .d1(q_23_11),
    .q(q_24_11)
  );
  

  flop_with_mux u_24_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_11),
    .d1(q_23_12),
    .q(q_24_12)
  );
  

  flop_with_mux u_24_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_12),
    .d1(q_23_13),
    .q(q_24_13)
  );
  

  flop_with_mux u_24_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_13),
    .d1(q_23_14),
    .q(q_24_14)
  );
  

  flop_with_mux u_24_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_14),
    .d1(q_23_15),
    .q(q_24_15)
  );
  

  flop_with_mux u_24_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_15),
    .d1(q_23_16),
    .q(q_24_16)
  );
  

  flop_with_mux u_24_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_16),
    .d1(q_23_17),
    .q(q_24_17)
  );
  

  flop_with_mux u_24_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_17),
    .d1(q_23_18),
    .q(q_24_18)
  );
  

  flop_with_mux u_24_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_18),
    .d1(q_23_19),
    .q(q_24_19)
  );
  

  flop_with_mux u_24_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_19),
    .d1(q_23_20),
    .q(q_24_20)
  );
  

  flop_with_mux u_24_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_20),
    .d1(q_23_21),
    .q(q_24_21)
  );
  

  flop_with_mux u_24_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_21),
    .d1(q_23_22),
    .q(q_24_22)
  );
  

  flop_with_mux u_24_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_22),
    .d1(q_23_23),
    .q(q_24_23)
  );
  

  flop_with_mux u_24_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_23),
    .d1(q_23_24),
    .q(q_24_24)
  );
  

  flop_with_mux u_24_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_24),
    .d1(q_23_25),
    .q(q_24_25)
  );
  

  flop_with_mux u_24_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_25),
    .d1(q_23_26),
    .q(q_24_26)
  );
  

  flop_with_mux u_24_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_26),
    .d1(q_23_27),
    .q(q_24_27)
  );
  

  flop_with_mux u_24_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_27),
    .d1(q_23_28),
    .q(q_24_28)
  );
  

  flop_with_mux u_24_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_28),
    .d1(q_23_29),
    .q(q_24_29)
  );
  

  flop_with_mux u_24_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_29),
    .d1(q_23_30),
    .q(q_24_30)
  );
  

  flop_with_mux u_24_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_30),
    .d1(q_23_31),
    .q(q_24_31)
  );
  

  flop_with_mux u_24_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_31),
    .d1(q_23_32),
    .q(q_24_32)
  );
  

  flop_with_mux u_24_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_32),
    .d1(q_23_33),
    .q(q_24_33)
  );
  

  flop_with_mux u_24_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_33),
    .d1(q_23_34),
    .q(q_24_34)
  );
  

  flop_with_mux u_24_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_34),
    .d1(q_23_35),
    .q(q_24_35)
  );
  

  flop_with_mux u_24_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_35),
    .d1(q_23_36),
    .q(q_24_36)
  );
  

  flop_with_mux u_24_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_36),
    .d1(q_23_37),
    .q(q_24_37)
  );
  

  flop_with_mux u_24_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_37),
    .d1(q_23_38),
    .q(q_24_38)
  );
  

  flop_with_mux u_24_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_24_38),
    .d1(q_23_39),
    .q(q_24_39)
  );
  

  flop_with_mux u_25_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_minus1),
    .d1(q_24_0),
    .q(q_25_0)
  );
  

  flop_with_mux u_25_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_0),
    .d1(q_24_1),
    .q(q_25_1)
  );
  

  flop_with_mux u_25_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_1),
    .d1(q_24_2),
    .q(q_25_2)
  );
  

  flop_with_mux u_25_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_2),
    .d1(q_24_3),
    .q(q_25_3)
  );
  

  flop_with_mux u_25_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_3),
    .d1(q_24_4),
    .q(q_25_4)
  );
  

  flop_with_mux u_25_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_4),
    .d1(q_24_5),
    .q(q_25_5)
  );
  

  flop_with_mux u_25_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_5),
    .d1(q_24_6),
    .q(q_25_6)
  );
  

  flop_with_mux u_25_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_6),
    .d1(q_24_7),
    .q(q_25_7)
  );
  

  flop_with_mux u_25_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_7),
    .d1(q_24_8),
    .q(q_25_8)
  );
  

  flop_with_mux u_25_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_8),
    .d1(q_24_9),
    .q(q_25_9)
  );
  

  flop_with_mux u_25_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_9),
    .d1(q_24_10),
    .q(q_25_10)
  );
  

  flop_with_mux u_25_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_10),
    .d1(q_24_11),
    .q(q_25_11)
  );
  

  flop_with_mux u_25_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_11),
    .d1(q_24_12),
    .q(q_25_12)
  );
  

  flop_with_mux u_25_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_12),
    .d1(q_24_13),
    .q(q_25_13)
  );
  

  flop_with_mux u_25_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_13),
    .d1(q_24_14),
    .q(q_25_14)
  );
  

  flop_with_mux u_25_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_14),
    .d1(q_24_15),
    .q(q_25_15)
  );
  

  flop_with_mux u_25_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_15),
    .d1(q_24_16),
    .q(q_25_16)
  );
  

  flop_with_mux u_25_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_16),
    .d1(q_24_17),
    .q(q_25_17)
  );
  

  flop_with_mux u_25_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_17),
    .d1(q_24_18),
    .q(q_25_18)
  );
  

  flop_with_mux u_25_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_18),
    .d1(q_24_19),
    .q(q_25_19)
  );
  

  flop_with_mux u_25_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_19),
    .d1(q_24_20),
    .q(q_25_20)
  );
  

  flop_with_mux u_25_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_20),
    .d1(q_24_21),
    .q(q_25_21)
  );
  

  flop_with_mux u_25_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_21),
    .d1(q_24_22),
    .q(q_25_22)
  );
  

  flop_with_mux u_25_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_22),
    .d1(q_24_23),
    .q(q_25_23)
  );
  

  flop_with_mux u_25_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_23),
    .d1(q_24_24),
    .q(q_25_24)
  );
  

  flop_with_mux u_25_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_24),
    .d1(q_24_25),
    .q(q_25_25)
  );
  

  flop_with_mux u_25_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_25),
    .d1(q_24_26),
    .q(q_25_26)
  );
  

  flop_with_mux u_25_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_26),
    .d1(q_24_27),
    .q(q_25_27)
  );
  

  flop_with_mux u_25_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_27),
    .d1(q_24_28),
    .q(q_25_28)
  );
  

  flop_with_mux u_25_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_28),
    .d1(q_24_29),
    .q(q_25_29)
  );
  

  flop_with_mux u_25_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_29),
    .d1(q_24_30),
    .q(q_25_30)
  );
  

  flop_with_mux u_25_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_30),
    .d1(q_24_31),
    .q(q_25_31)
  );
  

  flop_with_mux u_25_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_31),
    .d1(q_24_32),
    .q(q_25_32)
  );
  

  flop_with_mux u_25_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_32),
    .d1(q_24_33),
    .q(q_25_33)
  );
  

  flop_with_mux u_25_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_33),
    .d1(q_24_34),
    .q(q_25_34)
  );
  

  flop_with_mux u_25_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_34),
    .d1(q_24_35),
    .q(q_25_35)
  );
  

  flop_with_mux u_25_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_35),
    .d1(q_24_36),
    .q(q_25_36)
  );
  

  flop_with_mux u_25_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_36),
    .d1(q_24_37),
    .q(q_25_37)
  );
  

  flop_with_mux u_25_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_37),
    .d1(q_24_38),
    .q(q_25_38)
  );
  

  flop_with_mux u_25_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_25_38),
    .d1(q_24_39),
    .q(q_25_39)
  );
  

  flop_with_mux u_26_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_minus1),
    .d1(q_25_0),
    .q(q_26_0)
  );
  

  flop_with_mux u_26_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_0),
    .d1(q_25_1),
    .q(q_26_1)
  );
  

  flop_with_mux u_26_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_1),
    .d1(q_25_2),
    .q(q_26_2)
  );
  

  flop_with_mux u_26_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_2),
    .d1(q_25_3),
    .q(q_26_3)
  );
  

  flop_with_mux u_26_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_3),
    .d1(q_25_4),
    .q(q_26_4)
  );
  

  flop_with_mux u_26_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_4),
    .d1(q_25_5),
    .q(q_26_5)
  );
  

  flop_with_mux u_26_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_5),
    .d1(q_25_6),
    .q(q_26_6)
  );
  

  flop_with_mux u_26_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_6),
    .d1(q_25_7),
    .q(q_26_7)
  );
  

  flop_with_mux u_26_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_7),
    .d1(q_25_8),
    .q(q_26_8)
  );
  

  flop_with_mux u_26_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_8),
    .d1(q_25_9),
    .q(q_26_9)
  );
  

  flop_with_mux u_26_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_9),
    .d1(q_25_10),
    .q(q_26_10)
  );
  

  flop_with_mux u_26_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_10),
    .d1(q_25_11),
    .q(q_26_11)
  );
  

  flop_with_mux u_26_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_11),
    .d1(q_25_12),
    .q(q_26_12)
  );
  

  flop_with_mux u_26_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_12),
    .d1(q_25_13),
    .q(q_26_13)
  );
  

  flop_with_mux u_26_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_13),
    .d1(q_25_14),
    .q(q_26_14)
  );
  

  flop_with_mux u_26_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_14),
    .d1(q_25_15),
    .q(q_26_15)
  );
  

  flop_with_mux u_26_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_15),
    .d1(q_25_16),
    .q(q_26_16)
  );
  

  flop_with_mux u_26_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_16),
    .d1(q_25_17),
    .q(q_26_17)
  );
  

  flop_with_mux u_26_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_17),
    .d1(q_25_18),
    .q(q_26_18)
  );
  

  flop_with_mux u_26_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_18),
    .d1(q_25_19),
    .q(q_26_19)
  );
  

  flop_with_mux u_26_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_19),
    .d1(q_25_20),
    .q(q_26_20)
  );
  

  flop_with_mux u_26_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_20),
    .d1(q_25_21),
    .q(q_26_21)
  );
  

  flop_with_mux u_26_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_21),
    .d1(q_25_22),
    .q(q_26_22)
  );
  

  flop_with_mux u_26_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_22),
    .d1(q_25_23),
    .q(q_26_23)
  );
  

  flop_with_mux u_26_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_23),
    .d1(q_25_24),
    .q(q_26_24)
  );
  

  flop_with_mux u_26_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_24),
    .d1(q_25_25),
    .q(q_26_25)
  );
  

  flop_with_mux u_26_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_25),
    .d1(q_25_26),
    .q(q_26_26)
  );
  

  flop_with_mux u_26_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_26),
    .d1(q_25_27),
    .q(q_26_27)
  );
  

  flop_with_mux u_26_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_27),
    .d1(q_25_28),
    .q(q_26_28)
  );
  

  flop_with_mux u_26_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_28),
    .d1(q_25_29),
    .q(q_26_29)
  );
  

  flop_with_mux u_26_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_29),
    .d1(q_25_30),
    .q(q_26_30)
  );
  

  flop_with_mux u_26_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_30),
    .d1(q_25_31),
    .q(q_26_31)
  );
  

  flop_with_mux u_26_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_31),
    .d1(q_25_32),
    .q(q_26_32)
  );
  

  flop_with_mux u_26_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_32),
    .d1(q_25_33),
    .q(q_26_33)
  );
  

  flop_with_mux u_26_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_33),
    .d1(q_25_34),
    .q(q_26_34)
  );
  

  flop_with_mux u_26_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_34),
    .d1(q_25_35),
    .q(q_26_35)
  );
  

  flop_with_mux u_26_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_35),
    .d1(q_25_36),
    .q(q_26_36)
  );
  

  flop_with_mux u_26_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_36),
    .d1(q_25_37),
    .q(q_26_37)
  );
  

  flop_with_mux u_26_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_37),
    .d1(q_25_38),
    .q(q_26_38)
  );
  

  flop_with_mux u_26_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_26_38),
    .d1(q_25_39),
    .q(q_26_39)
  );
  

  flop_with_mux u_27_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_minus1),
    .d1(q_26_0),
    .q(q_27_0)
  );
  

  flop_with_mux u_27_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_0),
    .d1(q_26_1),
    .q(q_27_1)
  );
  

  flop_with_mux u_27_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_1),
    .d1(q_26_2),
    .q(q_27_2)
  );
  

  flop_with_mux u_27_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_2),
    .d1(q_26_3),
    .q(q_27_3)
  );
  

  flop_with_mux u_27_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_3),
    .d1(q_26_4),
    .q(q_27_4)
  );
  

  flop_with_mux u_27_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_4),
    .d1(q_26_5),
    .q(q_27_5)
  );
  

  flop_with_mux u_27_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_5),
    .d1(q_26_6),
    .q(q_27_6)
  );
  

  flop_with_mux u_27_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_6),
    .d1(q_26_7),
    .q(q_27_7)
  );
  

  flop_with_mux u_27_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_7),
    .d1(q_26_8),
    .q(q_27_8)
  );
  

  flop_with_mux u_27_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_8),
    .d1(q_26_9),
    .q(q_27_9)
  );
  

  flop_with_mux u_27_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_9),
    .d1(q_26_10),
    .q(q_27_10)
  );
  

  flop_with_mux u_27_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_10),
    .d1(q_26_11),
    .q(q_27_11)
  );
  

  flop_with_mux u_27_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_11),
    .d1(q_26_12),
    .q(q_27_12)
  );
  

  flop_with_mux u_27_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_12),
    .d1(q_26_13),
    .q(q_27_13)
  );
  

  flop_with_mux u_27_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_13),
    .d1(q_26_14),
    .q(q_27_14)
  );
  

  flop_with_mux u_27_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_14),
    .d1(q_26_15),
    .q(q_27_15)
  );
  

  flop_with_mux u_27_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_15),
    .d1(q_26_16),
    .q(q_27_16)
  );
  

  flop_with_mux u_27_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_16),
    .d1(q_26_17),
    .q(q_27_17)
  );
  

  flop_with_mux u_27_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_17),
    .d1(q_26_18),
    .q(q_27_18)
  );
  

  flop_with_mux u_27_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_18),
    .d1(q_26_19),
    .q(q_27_19)
  );
  

  flop_with_mux u_27_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_19),
    .d1(q_26_20),
    .q(q_27_20)
  );
  

  flop_with_mux u_27_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_20),
    .d1(q_26_21),
    .q(q_27_21)
  );
  

  flop_with_mux u_27_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_21),
    .d1(q_26_22),
    .q(q_27_22)
  );
  

  flop_with_mux u_27_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_22),
    .d1(q_26_23),
    .q(q_27_23)
  );
  

  flop_with_mux u_27_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_23),
    .d1(q_26_24),
    .q(q_27_24)
  );
  

  flop_with_mux u_27_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_24),
    .d1(q_26_25),
    .q(q_27_25)
  );
  

  flop_with_mux u_27_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_25),
    .d1(q_26_26),
    .q(q_27_26)
  );
  

  flop_with_mux u_27_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_26),
    .d1(q_26_27),
    .q(q_27_27)
  );
  

  flop_with_mux u_27_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_27),
    .d1(q_26_28),
    .q(q_27_28)
  );
  

  flop_with_mux u_27_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_28),
    .d1(q_26_29),
    .q(q_27_29)
  );
  

  flop_with_mux u_27_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_29),
    .d1(q_26_30),
    .q(q_27_30)
  );
  

  flop_with_mux u_27_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_30),
    .d1(q_26_31),
    .q(q_27_31)
  );
  

  flop_with_mux u_27_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_31),
    .d1(q_26_32),
    .q(q_27_32)
  );
  

  flop_with_mux u_27_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_32),
    .d1(q_26_33),
    .q(q_27_33)
  );
  

  flop_with_mux u_27_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_33),
    .d1(q_26_34),
    .q(q_27_34)
  );
  

  flop_with_mux u_27_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_34),
    .d1(q_26_35),
    .q(q_27_35)
  );
  

  flop_with_mux u_27_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_35),
    .d1(q_26_36),
    .q(q_27_36)
  );
  

  flop_with_mux u_27_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_36),
    .d1(q_26_37),
    .q(q_27_37)
  );
  

  flop_with_mux u_27_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_37),
    .d1(q_26_38),
    .q(q_27_38)
  );
  

  flop_with_mux u_27_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_27_38),
    .d1(q_26_39),
    .q(q_27_39)
  );
  

  flop_with_mux u_28_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_minus1),
    .d1(q_27_0),
    .q(q_28_0)
  );
  

  flop_with_mux u_28_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_0),
    .d1(q_27_1),
    .q(q_28_1)
  );
  

  flop_with_mux u_28_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_1),
    .d1(q_27_2),
    .q(q_28_2)
  );
  

  flop_with_mux u_28_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_2),
    .d1(q_27_3),
    .q(q_28_3)
  );
  

  flop_with_mux u_28_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_3),
    .d1(q_27_4),
    .q(q_28_4)
  );
  

  flop_with_mux u_28_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_4),
    .d1(q_27_5),
    .q(q_28_5)
  );
  

  flop_with_mux u_28_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_5),
    .d1(q_27_6),
    .q(q_28_6)
  );
  

  flop_with_mux u_28_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_6),
    .d1(q_27_7),
    .q(q_28_7)
  );
  

  flop_with_mux u_28_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_7),
    .d1(q_27_8),
    .q(q_28_8)
  );
  

  flop_with_mux u_28_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_8),
    .d1(q_27_9),
    .q(q_28_9)
  );
  

  flop_with_mux u_28_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_9),
    .d1(q_27_10),
    .q(q_28_10)
  );
  

  flop_with_mux u_28_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_10),
    .d1(q_27_11),
    .q(q_28_11)
  );
  

  flop_with_mux u_28_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_11),
    .d1(q_27_12),
    .q(q_28_12)
  );
  

  flop_with_mux u_28_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_12),
    .d1(q_27_13),
    .q(q_28_13)
  );
  

  flop_with_mux u_28_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_13),
    .d1(q_27_14),
    .q(q_28_14)
  );
  

  flop_with_mux u_28_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_14),
    .d1(q_27_15),
    .q(q_28_15)
  );
  

  flop_with_mux u_28_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_15),
    .d1(q_27_16),
    .q(q_28_16)
  );
  

  flop_with_mux u_28_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_16),
    .d1(q_27_17),
    .q(q_28_17)
  );
  

  flop_with_mux u_28_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_17),
    .d1(q_27_18),
    .q(q_28_18)
  );
  

  flop_with_mux u_28_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_18),
    .d1(q_27_19),
    .q(q_28_19)
  );
  

  flop_with_mux u_28_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_19),
    .d1(q_27_20),
    .q(q_28_20)
  );
  

  flop_with_mux u_28_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_20),
    .d1(q_27_21),
    .q(q_28_21)
  );
  

  flop_with_mux u_28_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_21),
    .d1(q_27_22),
    .q(q_28_22)
  );
  

  flop_with_mux u_28_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_22),
    .d1(q_27_23),
    .q(q_28_23)
  );
  

  flop_with_mux u_28_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_23),
    .d1(q_27_24),
    .q(q_28_24)
  );
  

  flop_with_mux u_28_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_24),
    .d1(q_27_25),
    .q(q_28_25)
  );
  

  flop_with_mux u_28_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_25),
    .d1(q_27_26),
    .q(q_28_26)
  );
  

  flop_with_mux u_28_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_26),
    .d1(q_27_27),
    .q(q_28_27)
  );
  

  flop_with_mux u_28_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_27),
    .d1(q_27_28),
    .q(q_28_28)
  );
  

  flop_with_mux u_28_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_28),
    .d1(q_27_29),
    .q(q_28_29)
  );
  

  flop_with_mux u_28_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_29),
    .d1(q_27_30),
    .q(q_28_30)
  );
  

  flop_with_mux u_28_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_30),
    .d1(q_27_31),
    .q(q_28_31)
  );
  

  flop_with_mux u_28_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_31),
    .d1(q_27_32),
    .q(q_28_32)
  );
  

  flop_with_mux u_28_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_32),
    .d1(q_27_33),
    .q(q_28_33)
  );
  

  flop_with_mux u_28_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_33),
    .d1(q_27_34),
    .q(q_28_34)
  );
  

  flop_with_mux u_28_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_34),
    .d1(q_27_35),
    .q(q_28_35)
  );
  

  flop_with_mux u_28_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_35),
    .d1(q_27_36),
    .q(q_28_36)
  );
  

  flop_with_mux u_28_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_36),
    .d1(q_27_37),
    .q(q_28_37)
  );
  

  flop_with_mux u_28_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_37),
    .d1(q_27_38),
    .q(q_28_38)
  );
  

  flop_with_mux u_28_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_28_38),
    .d1(q_27_39),
    .q(q_28_39)
  );
  

  flop_with_mux u_29_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_minus1),
    .d1(q_28_0),
    .q(q_29_0)
  );
  

  flop_with_mux u_29_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_0),
    .d1(q_28_1),
    .q(q_29_1)
  );
  

  flop_with_mux u_29_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_1),
    .d1(q_28_2),
    .q(q_29_2)
  );
  

  flop_with_mux u_29_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_2),
    .d1(q_28_3),
    .q(q_29_3)
  );
  

  flop_with_mux u_29_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_3),
    .d1(q_28_4),
    .q(q_29_4)
  );
  

  flop_with_mux u_29_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_4),
    .d1(q_28_5),
    .q(q_29_5)
  );
  

  flop_with_mux u_29_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_5),
    .d1(q_28_6),
    .q(q_29_6)
  );
  

  flop_with_mux u_29_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_6),
    .d1(q_28_7),
    .q(q_29_7)
  );
  

  flop_with_mux u_29_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_7),
    .d1(q_28_8),
    .q(q_29_8)
  );
  

  flop_with_mux u_29_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_8),
    .d1(q_28_9),
    .q(q_29_9)
  );
  

  flop_with_mux u_29_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_9),
    .d1(q_28_10),
    .q(q_29_10)
  );
  

  flop_with_mux u_29_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_10),
    .d1(q_28_11),
    .q(q_29_11)
  );
  

  flop_with_mux u_29_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_11),
    .d1(q_28_12),
    .q(q_29_12)
  );
  

  flop_with_mux u_29_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_12),
    .d1(q_28_13),
    .q(q_29_13)
  );
  

  flop_with_mux u_29_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_13),
    .d1(q_28_14),
    .q(q_29_14)
  );
  

  flop_with_mux u_29_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_14),
    .d1(q_28_15),
    .q(q_29_15)
  );
  

  flop_with_mux u_29_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_15),
    .d1(q_28_16),
    .q(q_29_16)
  );
  

  flop_with_mux u_29_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_16),
    .d1(q_28_17),
    .q(q_29_17)
  );
  

  flop_with_mux u_29_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_17),
    .d1(q_28_18),
    .q(q_29_18)
  );
  

  flop_with_mux u_29_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_18),
    .d1(q_28_19),
    .q(q_29_19)
  );
  

  flop_with_mux u_29_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_19),
    .d1(q_28_20),
    .q(q_29_20)
  );
  

  flop_with_mux u_29_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_20),
    .d1(q_28_21),
    .q(q_29_21)
  );
  

  flop_with_mux u_29_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_21),
    .d1(q_28_22),
    .q(q_29_22)
  );
  

  flop_with_mux u_29_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_22),
    .d1(q_28_23),
    .q(q_29_23)
  );
  

  flop_with_mux u_29_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_23),
    .d1(q_28_24),
    .q(q_29_24)
  );
  

  flop_with_mux u_29_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_24),
    .d1(q_28_25),
    .q(q_29_25)
  );
  

  flop_with_mux u_29_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_25),
    .d1(q_28_26),
    .q(q_29_26)
  );
  

  flop_with_mux u_29_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_26),
    .d1(q_28_27),
    .q(q_29_27)
  );
  

  flop_with_mux u_29_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_27),
    .d1(q_28_28),
    .q(q_29_28)
  );
  

  flop_with_mux u_29_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_28),
    .d1(q_28_29),
    .q(q_29_29)
  );
  

  flop_with_mux u_29_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_29),
    .d1(q_28_30),
    .q(q_29_30)
  );
  

  flop_with_mux u_29_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_30),
    .d1(q_28_31),
    .q(q_29_31)
  );
  

  flop_with_mux u_29_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_31),
    .d1(q_28_32),
    .q(q_29_32)
  );
  

  flop_with_mux u_29_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_32),
    .d1(q_28_33),
    .q(q_29_33)
  );
  

  flop_with_mux u_29_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_33),
    .d1(q_28_34),
    .q(q_29_34)
  );
  

  flop_with_mux u_29_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_34),
    .d1(q_28_35),
    .q(q_29_35)
  );
  

  flop_with_mux u_29_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_35),
    .d1(q_28_36),
    .q(q_29_36)
  );
  

  flop_with_mux u_29_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_36),
    .d1(q_28_37),
    .q(q_29_37)
  );
  

  flop_with_mux u_29_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_37),
    .d1(q_28_38),
    .q(q_29_38)
  );
  

  flop_with_mux u_29_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_29_38),
    .d1(q_28_39),
    .q(q_29_39)
  );
  

  flop_with_mux u_30_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_minus1),
    .d1(q_29_0),
    .q(q_30_0)
  );
  

  flop_with_mux u_30_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_0),
    .d1(q_29_1),
    .q(q_30_1)
  );
  

  flop_with_mux u_30_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_1),
    .d1(q_29_2),
    .q(q_30_2)
  );
  

  flop_with_mux u_30_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_2),
    .d1(q_29_3),
    .q(q_30_3)
  );
  

  flop_with_mux u_30_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_3),
    .d1(q_29_4),
    .q(q_30_4)
  );
  

  flop_with_mux u_30_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_4),
    .d1(q_29_5),
    .q(q_30_5)
  );
  

  flop_with_mux u_30_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_5),
    .d1(q_29_6),
    .q(q_30_6)
  );
  

  flop_with_mux u_30_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_6),
    .d1(q_29_7),
    .q(q_30_7)
  );
  

  flop_with_mux u_30_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_7),
    .d1(q_29_8),
    .q(q_30_8)
  );
  

  flop_with_mux u_30_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_8),
    .d1(q_29_9),
    .q(q_30_9)
  );
  

  flop_with_mux u_30_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_9),
    .d1(q_29_10),
    .q(q_30_10)
  );
  

  flop_with_mux u_30_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_10),
    .d1(q_29_11),
    .q(q_30_11)
  );
  

  flop_with_mux u_30_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_11),
    .d1(q_29_12),
    .q(q_30_12)
  );
  

  flop_with_mux u_30_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_12),
    .d1(q_29_13),
    .q(q_30_13)
  );
  

  flop_with_mux u_30_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_13),
    .d1(q_29_14),
    .q(q_30_14)
  );
  

  flop_with_mux u_30_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_14),
    .d1(q_29_15),
    .q(q_30_15)
  );
  

  flop_with_mux u_30_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_15),
    .d1(q_29_16),
    .q(q_30_16)
  );
  

  flop_with_mux u_30_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_16),
    .d1(q_29_17),
    .q(q_30_17)
  );
  

  flop_with_mux u_30_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_17),
    .d1(q_29_18),
    .q(q_30_18)
  );
  

  flop_with_mux u_30_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_18),
    .d1(q_29_19),
    .q(q_30_19)
  );
  

  flop_with_mux u_30_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_19),
    .d1(q_29_20),
    .q(q_30_20)
  );
  

  flop_with_mux u_30_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_20),
    .d1(q_29_21),
    .q(q_30_21)
  );
  

  flop_with_mux u_30_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_21),
    .d1(q_29_22),
    .q(q_30_22)
  );
  

  flop_with_mux u_30_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_22),
    .d1(q_29_23),
    .q(q_30_23)
  );
  

  flop_with_mux u_30_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_23),
    .d1(q_29_24),
    .q(q_30_24)
  );
  

  flop_with_mux u_30_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_24),
    .d1(q_29_25),
    .q(q_30_25)
  );
  

  flop_with_mux u_30_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_25),
    .d1(q_29_26),
    .q(q_30_26)
  );
  

  flop_with_mux u_30_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_26),
    .d1(q_29_27),
    .q(q_30_27)
  );
  

  flop_with_mux u_30_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_27),
    .d1(q_29_28),
    .q(q_30_28)
  );
  

  flop_with_mux u_30_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_28),
    .d1(q_29_29),
    .q(q_30_29)
  );
  

  flop_with_mux u_30_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_29),
    .d1(q_29_30),
    .q(q_30_30)
  );
  

  flop_with_mux u_30_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_30),
    .d1(q_29_31),
    .q(q_30_31)
  );
  

  flop_with_mux u_30_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_31),
    .d1(q_29_32),
    .q(q_30_32)
  );
  

  flop_with_mux u_30_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_32),
    .d1(q_29_33),
    .q(q_30_33)
  );
  

  flop_with_mux u_30_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_33),
    .d1(q_29_34),
    .q(q_30_34)
  );
  

  flop_with_mux u_30_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_34),
    .d1(q_29_35),
    .q(q_30_35)
  );
  

  flop_with_mux u_30_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_35),
    .d1(q_29_36),
    .q(q_30_36)
  );
  

  flop_with_mux u_30_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_36),
    .d1(q_29_37),
    .q(q_30_37)
  );
  

  flop_with_mux u_30_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_37),
    .d1(q_29_38),
    .q(q_30_38)
  );
  

  flop_with_mux u_30_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_30_38),
    .d1(q_29_39),
    .q(q_30_39)
  );
  

  flop_with_mux u_31_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_minus1),
    .d1(q_30_0),
    .q(q_31_0)
  );
  

  flop_with_mux u_31_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_0),
    .d1(q_30_1),
    .q(q_31_1)
  );
  

  flop_with_mux u_31_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_1),
    .d1(q_30_2),
    .q(q_31_2)
  );
  

  flop_with_mux u_31_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_2),
    .d1(q_30_3),
    .q(q_31_3)
  );
  

  flop_with_mux u_31_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_3),
    .d1(q_30_4),
    .q(q_31_4)
  );
  

  flop_with_mux u_31_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_4),
    .d1(q_30_5),
    .q(q_31_5)
  );
  

  flop_with_mux u_31_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_5),
    .d1(q_30_6),
    .q(q_31_6)
  );
  

  flop_with_mux u_31_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_6),
    .d1(q_30_7),
    .q(q_31_7)
  );
  

  flop_with_mux u_31_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_7),
    .d1(q_30_8),
    .q(q_31_8)
  );
  

  flop_with_mux u_31_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_8),
    .d1(q_30_9),
    .q(q_31_9)
  );
  

  flop_with_mux u_31_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_9),
    .d1(q_30_10),
    .q(q_31_10)
  );
  

  flop_with_mux u_31_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_10),
    .d1(q_30_11),
    .q(q_31_11)
  );
  

  flop_with_mux u_31_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_11),
    .d1(q_30_12),
    .q(q_31_12)
  );
  

  flop_with_mux u_31_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_12),
    .d1(q_30_13),
    .q(q_31_13)
  );
  

  flop_with_mux u_31_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_13),
    .d1(q_30_14),
    .q(q_31_14)
  );
  

  flop_with_mux u_31_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_14),
    .d1(q_30_15),
    .q(q_31_15)
  );
  

  flop_with_mux u_31_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_15),
    .d1(q_30_16),
    .q(q_31_16)
  );
  

  flop_with_mux u_31_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_16),
    .d1(q_30_17),
    .q(q_31_17)
  );
  

  flop_with_mux u_31_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_17),
    .d1(q_30_18),
    .q(q_31_18)
  );
  

  flop_with_mux u_31_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_18),
    .d1(q_30_19),
    .q(q_31_19)
  );
  

  flop_with_mux u_31_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_19),
    .d1(q_30_20),
    .q(q_31_20)
  );
  

  flop_with_mux u_31_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_20),
    .d1(q_30_21),
    .q(q_31_21)
  );
  

  flop_with_mux u_31_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_21),
    .d1(q_30_22),
    .q(q_31_22)
  );
  

  flop_with_mux u_31_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_22),
    .d1(q_30_23),
    .q(q_31_23)
  );
  

  flop_with_mux u_31_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_23),
    .d1(q_30_24),
    .q(q_31_24)
  );
  

  flop_with_mux u_31_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_24),
    .d1(q_30_25),
    .q(q_31_25)
  );
  

  flop_with_mux u_31_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_25),
    .d1(q_30_26),
    .q(q_31_26)
  );
  

  flop_with_mux u_31_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_26),
    .d1(q_30_27),
    .q(q_31_27)
  );
  

  flop_with_mux u_31_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_27),
    .d1(q_30_28),
    .q(q_31_28)
  );
  

  flop_with_mux u_31_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_28),
    .d1(q_30_29),
    .q(q_31_29)
  );
  

  flop_with_mux u_31_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_29),
    .d1(q_30_30),
    .q(q_31_30)
  );
  

  flop_with_mux u_31_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_30),
    .d1(q_30_31),
    .q(q_31_31)
  );
  

  flop_with_mux u_31_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_31),
    .d1(q_30_32),
    .q(q_31_32)
  );
  

  flop_with_mux u_31_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_32),
    .d1(q_30_33),
    .q(q_31_33)
  );
  

  flop_with_mux u_31_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_33),
    .d1(q_30_34),
    .q(q_31_34)
  );
  

  flop_with_mux u_31_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_34),
    .d1(q_30_35),
    .q(q_31_35)
  );
  

  flop_with_mux u_31_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_35),
    .d1(q_30_36),
    .q(q_31_36)
  );
  

  flop_with_mux u_31_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_36),
    .d1(q_30_37),
    .q(q_31_37)
  );
  

  flop_with_mux u_31_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_37),
    .d1(q_30_38),
    .q(q_31_38)
  );
  

  flop_with_mux u_31_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_31_38),
    .d1(q_30_39),
    .q(q_31_39)
  );
  

  flop_with_mux u_32_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_minus1),
    .d1(q_31_0),
    .q(q_32_0)
  );
  

  flop_with_mux u_32_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_0),
    .d1(q_31_1),
    .q(q_32_1)
  );
  

  flop_with_mux u_32_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_1),
    .d1(q_31_2),
    .q(q_32_2)
  );
  

  flop_with_mux u_32_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_2),
    .d1(q_31_3),
    .q(q_32_3)
  );
  

  flop_with_mux u_32_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_3),
    .d1(q_31_4),
    .q(q_32_4)
  );
  

  flop_with_mux u_32_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_4),
    .d1(q_31_5),
    .q(q_32_5)
  );
  

  flop_with_mux u_32_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_5),
    .d1(q_31_6),
    .q(q_32_6)
  );
  

  flop_with_mux u_32_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_6),
    .d1(q_31_7),
    .q(q_32_7)
  );
  

  flop_with_mux u_32_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_7),
    .d1(q_31_8),
    .q(q_32_8)
  );
  

  flop_with_mux u_32_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_8),
    .d1(q_31_9),
    .q(q_32_9)
  );
  

  flop_with_mux u_32_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_9),
    .d1(q_31_10),
    .q(q_32_10)
  );
  

  flop_with_mux u_32_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_10),
    .d1(q_31_11),
    .q(q_32_11)
  );
  

  flop_with_mux u_32_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_11),
    .d1(q_31_12),
    .q(q_32_12)
  );
  

  flop_with_mux u_32_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_12),
    .d1(q_31_13),
    .q(q_32_13)
  );
  

  flop_with_mux u_32_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_13),
    .d1(q_31_14),
    .q(q_32_14)
  );
  

  flop_with_mux u_32_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_14),
    .d1(q_31_15),
    .q(q_32_15)
  );
  

  flop_with_mux u_32_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_15),
    .d1(q_31_16),
    .q(q_32_16)
  );
  

  flop_with_mux u_32_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_16),
    .d1(q_31_17),
    .q(q_32_17)
  );
  

  flop_with_mux u_32_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_17),
    .d1(q_31_18),
    .q(q_32_18)
  );
  

  flop_with_mux u_32_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_18),
    .d1(q_31_19),
    .q(q_32_19)
  );
  

  flop_with_mux u_32_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_19),
    .d1(q_31_20),
    .q(q_32_20)
  );
  

  flop_with_mux u_32_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_20),
    .d1(q_31_21),
    .q(q_32_21)
  );
  

  flop_with_mux u_32_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_21),
    .d1(q_31_22),
    .q(q_32_22)
  );
  

  flop_with_mux u_32_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_22),
    .d1(q_31_23),
    .q(q_32_23)
  );
  

  flop_with_mux u_32_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_23),
    .d1(q_31_24),
    .q(q_32_24)
  );
  

  flop_with_mux u_32_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_24),
    .d1(q_31_25),
    .q(q_32_25)
  );
  

  flop_with_mux u_32_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_25),
    .d1(q_31_26),
    .q(q_32_26)
  );
  

  flop_with_mux u_32_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_26),
    .d1(q_31_27),
    .q(q_32_27)
  );
  

  flop_with_mux u_32_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_27),
    .d1(q_31_28),
    .q(q_32_28)
  );
  

  flop_with_mux u_32_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_28),
    .d1(q_31_29),
    .q(q_32_29)
  );
  

  flop_with_mux u_32_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_29),
    .d1(q_31_30),
    .q(q_32_30)
  );
  

  flop_with_mux u_32_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_30),
    .d1(q_31_31),
    .q(q_32_31)
  );
  

  flop_with_mux u_32_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_31),
    .d1(q_31_32),
    .q(q_32_32)
  );
  

  flop_with_mux u_32_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_32),
    .d1(q_31_33),
    .q(q_32_33)
  );
  

  flop_with_mux u_32_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_33),
    .d1(q_31_34),
    .q(q_32_34)
  );
  

  flop_with_mux u_32_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_34),
    .d1(q_31_35),
    .q(q_32_35)
  );
  

  flop_with_mux u_32_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_35),
    .d1(q_31_36),
    .q(q_32_36)
  );
  

  flop_with_mux u_32_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_36),
    .d1(q_31_37),
    .q(q_32_37)
  );
  

  flop_with_mux u_32_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_37),
    .d1(q_31_38),
    .q(q_32_38)
  );
  

  flop_with_mux u_32_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_32_38),
    .d1(q_31_39),
    .q(q_32_39)
  );
  

  flop_with_mux u_33_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_minus1),
    .d1(q_32_0),
    .q(q_33_0)
  );
  

  flop_with_mux u_33_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_0),
    .d1(q_32_1),
    .q(q_33_1)
  );
  

  flop_with_mux u_33_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_1),
    .d1(q_32_2),
    .q(q_33_2)
  );
  

  flop_with_mux u_33_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_2),
    .d1(q_32_3),
    .q(q_33_3)
  );
  

  flop_with_mux u_33_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_3),
    .d1(q_32_4),
    .q(q_33_4)
  );
  

  flop_with_mux u_33_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_4),
    .d1(q_32_5),
    .q(q_33_5)
  );
  

  flop_with_mux u_33_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_5),
    .d1(q_32_6),
    .q(q_33_6)
  );
  

  flop_with_mux u_33_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_6),
    .d1(q_32_7),
    .q(q_33_7)
  );
  

  flop_with_mux u_33_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_7),
    .d1(q_32_8),
    .q(q_33_8)
  );
  

  flop_with_mux u_33_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_8),
    .d1(q_32_9),
    .q(q_33_9)
  );
  

  flop_with_mux u_33_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_9),
    .d1(q_32_10),
    .q(q_33_10)
  );
  

  flop_with_mux u_33_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_10),
    .d1(q_32_11),
    .q(q_33_11)
  );
  

  flop_with_mux u_33_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_11),
    .d1(q_32_12),
    .q(q_33_12)
  );
  

  flop_with_mux u_33_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_12),
    .d1(q_32_13),
    .q(q_33_13)
  );
  

  flop_with_mux u_33_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_13),
    .d1(q_32_14),
    .q(q_33_14)
  );
  

  flop_with_mux u_33_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_14),
    .d1(q_32_15),
    .q(q_33_15)
  );
  

  flop_with_mux u_33_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_15),
    .d1(q_32_16),
    .q(q_33_16)
  );
  

  flop_with_mux u_33_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_16),
    .d1(q_32_17),
    .q(q_33_17)
  );
  

  flop_with_mux u_33_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_17),
    .d1(q_32_18),
    .q(q_33_18)
  );
  

  flop_with_mux u_33_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_18),
    .d1(q_32_19),
    .q(q_33_19)
  );
  

  flop_with_mux u_33_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_19),
    .d1(q_32_20),
    .q(q_33_20)
  );
  

  flop_with_mux u_33_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_20),
    .d1(q_32_21),
    .q(q_33_21)
  );
  

  flop_with_mux u_33_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_21),
    .d1(q_32_22),
    .q(q_33_22)
  );
  

  flop_with_mux u_33_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_22),
    .d1(q_32_23),
    .q(q_33_23)
  );
  

  flop_with_mux u_33_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_23),
    .d1(q_32_24),
    .q(q_33_24)
  );
  

  flop_with_mux u_33_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_24),
    .d1(q_32_25),
    .q(q_33_25)
  );
  

  flop_with_mux u_33_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_25),
    .d1(q_32_26),
    .q(q_33_26)
  );
  

  flop_with_mux u_33_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_26),
    .d1(q_32_27),
    .q(q_33_27)
  );
  

  flop_with_mux u_33_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_27),
    .d1(q_32_28),
    .q(q_33_28)
  );
  

  flop_with_mux u_33_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_28),
    .d1(q_32_29),
    .q(q_33_29)
  );
  

  flop_with_mux u_33_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_29),
    .d1(q_32_30),
    .q(q_33_30)
  );
  

  flop_with_mux u_33_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_30),
    .d1(q_32_31),
    .q(q_33_31)
  );
  

  flop_with_mux u_33_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_31),
    .d1(q_32_32),
    .q(q_33_32)
  );
  

  flop_with_mux u_33_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_32),
    .d1(q_32_33),
    .q(q_33_33)
  );
  

  flop_with_mux u_33_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_33),
    .d1(q_32_34),
    .q(q_33_34)
  );
  

  flop_with_mux u_33_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_34),
    .d1(q_32_35),
    .q(q_33_35)
  );
  

  flop_with_mux u_33_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_35),
    .d1(q_32_36),
    .q(q_33_36)
  );
  

  flop_with_mux u_33_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_36),
    .d1(q_32_37),
    .q(q_33_37)
  );
  

  flop_with_mux u_33_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_37),
    .d1(q_32_38),
    .q(q_33_38)
  );
  

  flop_with_mux u_33_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_33_38),
    .d1(q_32_39),
    .q(q_33_39)
  );
  

  flop_with_mux u_34_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_minus1),
    .d1(q_33_0),
    .q(q_34_0)
  );
  

  flop_with_mux u_34_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_0),
    .d1(q_33_1),
    .q(q_34_1)
  );
  

  flop_with_mux u_34_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_1),
    .d1(q_33_2),
    .q(q_34_2)
  );
  

  flop_with_mux u_34_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_2),
    .d1(q_33_3),
    .q(q_34_3)
  );
  

  flop_with_mux u_34_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_3),
    .d1(q_33_4),
    .q(q_34_4)
  );
  

  flop_with_mux u_34_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_4),
    .d1(q_33_5),
    .q(q_34_5)
  );
  

  flop_with_mux u_34_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_5),
    .d1(q_33_6),
    .q(q_34_6)
  );
  

  flop_with_mux u_34_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_6),
    .d1(q_33_7),
    .q(q_34_7)
  );
  

  flop_with_mux u_34_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_7),
    .d1(q_33_8),
    .q(q_34_8)
  );
  

  flop_with_mux u_34_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_8),
    .d1(q_33_9),
    .q(q_34_9)
  );
  

  flop_with_mux u_34_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_9),
    .d1(q_33_10),
    .q(q_34_10)
  );
  

  flop_with_mux u_34_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_10),
    .d1(q_33_11),
    .q(q_34_11)
  );
  

  flop_with_mux u_34_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_11),
    .d1(q_33_12),
    .q(q_34_12)
  );
  

  flop_with_mux u_34_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_12),
    .d1(q_33_13),
    .q(q_34_13)
  );
  

  flop_with_mux u_34_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_13),
    .d1(q_33_14),
    .q(q_34_14)
  );
  

  flop_with_mux u_34_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_14),
    .d1(q_33_15),
    .q(q_34_15)
  );
  

  flop_with_mux u_34_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_15),
    .d1(q_33_16),
    .q(q_34_16)
  );
  

  flop_with_mux u_34_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_16),
    .d1(q_33_17),
    .q(q_34_17)
  );
  

  flop_with_mux u_34_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_17),
    .d1(q_33_18),
    .q(q_34_18)
  );
  

  flop_with_mux u_34_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_18),
    .d1(q_33_19),
    .q(q_34_19)
  );
  

  flop_with_mux u_34_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_19),
    .d1(q_33_20),
    .q(q_34_20)
  );
  

  flop_with_mux u_34_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_20),
    .d1(q_33_21),
    .q(q_34_21)
  );
  

  flop_with_mux u_34_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_21),
    .d1(q_33_22),
    .q(q_34_22)
  );
  

  flop_with_mux u_34_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_22),
    .d1(q_33_23),
    .q(q_34_23)
  );
  

  flop_with_mux u_34_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_23),
    .d1(q_33_24),
    .q(q_34_24)
  );
  

  flop_with_mux u_34_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_24),
    .d1(q_33_25),
    .q(q_34_25)
  );
  

  flop_with_mux u_34_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_25),
    .d1(q_33_26),
    .q(q_34_26)
  );
  

  flop_with_mux u_34_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_26),
    .d1(q_33_27),
    .q(q_34_27)
  );
  

  flop_with_mux u_34_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_27),
    .d1(q_33_28),
    .q(q_34_28)
  );
  

  flop_with_mux u_34_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_28),
    .d1(q_33_29),
    .q(q_34_29)
  );
  

  flop_with_mux u_34_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_29),
    .d1(q_33_30),
    .q(q_34_30)
  );
  

  flop_with_mux u_34_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_30),
    .d1(q_33_31),
    .q(q_34_31)
  );
  

  flop_with_mux u_34_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_31),
    .d1(q_33_32),
    .q(q_34_32)
  );
  

  flop_with_mux u_34_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_32),
    .d1(q_33_33),
    .q(q_34_33)
  );
  

  flop_with_mux u_34_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_33),
    .d1(q_33_34),
    .q(q_34_34)
  );
  

  flop_with_mux u_34_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_34),
    .d1(q_33_35),
    .q(q_34_35)
  );
  

  flop_with_mux u_34_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_35),
    .d1(q_33_36),
    .q(q_34_36)
  );
  

  flop_with_mux u_34_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_36),
    .d1(q_33_37),
    .q(q_34_37)
  );
  

  flop_with_mux u_34_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_37),
    .d1(q_33_38),
    .q(q_34_38)
  );
  

  flop_with_mux u_34_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_34_38),
    .d1(q_33_39),
    .q(q_34_39)
  );
  

  flop_with_mux u_35_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_minus1),
    .d1(q_34_0),
    .q(q_35_0)
  );
  

  flop_with_mux u_35_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_0),
    .d1(q_34_1),
    .q(q_35_1)
  );
  

  flop_with_mux u_35_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_1),
    .d1(q_34_2),
    .q(q_35_2)
  );
  

  flop_with_mux u_35_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_2),
    .d1(q_34_3),
    .q(q_35_3)
  );
  

  flop_with_mux u_35_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_3),
    .d1(q_34_4),
    .q(q_35_4)
  );
  

  flop_with_mux u_35_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_4),
    .d1(q_34_5),
    .q(q_35_5)
  );
  

  flop_with_mux u_35_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_5),
    .d1(q_34_6),
    .q(q_35_6)
  );
  

  flop_with_mux u_35_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_6),
    .d1(q_34_7),
    .q(q_35_7)
  );
  

  flop_with_mux u_35_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_7),
    .d1(q_34_8),
    .q(q_35_8)
  );
  

  flop_with_mux u_35_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_8),
    .d1(q_34_9),
    .q(q_35_9)
  );
  

  flop_with_mux u_35_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_9),
    .d1(q_34_10),
    .q(q_35_10)
  );
  

  flop_with_mux u_35_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_10),
    .d1(q_34_11),
    .q(q_35_11)
  );
  

  flop_with_mux u_35_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_11),
    .d1(q_34_12),
    .q(q_35_12)
  );
  

  flop_with_mux u_35_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_12),
    .d1(q_34_13),
    .q(q_35_13)
  );
  

  flop_with_mux u_35_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_13),
    .d1(q_34_14),
    .q(q_35_14)
  );
  

  flop_with_mux u_35_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_14),
    .d1(q_34_15),
    .q(q_35_15)
  );
  

  flop_with_mux u_35_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_15),
    .d1(q_34_16),
    .q(q_35_16)
  );
  

  flop_with_mux u_35_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_16),
    .d1(q_34_17),
    .q(q_35_17)
  );
  

  flop_with_mux u_35_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_17),
    .d1(q_34_18),
    .q(q_35_18)
  );
  

  flop_with_mux u_35_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_18),
    .d1(q_34_19),
    .q(q_35_19)
  );
  

  flop_with_mux u_35_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_19),
    .d1(q_34_20),
    .q(q_35_20)
  );
  

  flop_with_mux u_35_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_20),
    .d1(q_34_21),
    .q(q_35_21)
  );
  

  flop_with_mux u_35_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_21),
    .d1(q_34_22),
    .q(q_35_22)
  );
  

  flop_with_mux u_35_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_22),
    .d1(q_34_23),
    .q(q_35_23)
  );
  

  flop_with_mux u_35_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_23),
    .d1(q_34_24),
    .q(q_35_24)
  );
  

  flop_with_mux u_35_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_24),
    .d1(q_34_25),
    .q(q_35_25)
  );
  

  flop_with_mux u_35_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_25),
    .d1(q_34_26),
    .q(q_35_26)
  );
  

  flop_with_mux u_35_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_26),
    .d1(q_34_27),
    .q(q_35_27)
  );
  

  flop_with_mux u_35_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_27),
    .d1(q_34_28),
    .q(q_35_28)
  );
  

  flop_with_mux u_35_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_28),
    .d1(q_34_29),
    .q(q_35_29)
  );
  

  flop_with_mux u_35_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_29),
    .d1(q_34_30),
    .q(q_35_30)
  );
  

  flop_with_mux u_35_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_30),
    .d1(q_34_31),
    .q(q_35_31)
  );
  

  flop_with_mux u_35_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_31),
    .d1(q_34_32),
    .q(q_35_32)
  );
  

  flop_with_mux u_35_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_32),
    .d1(q_34_33),
    .q(q_35_33)
  );
  

  flop_with_mux u_35_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_33),
    .d1(q_34_34),
    .q(q_35_34)
  );
  

  flop_with_mux u_35_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_34),
    .d1(q_34_35),
    .q(q_35_35)
  );
  

  flop_with_mux u_35_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_35),
    .d1(q_34_36),
    .q(q_35_36)
  );
  

  flop_with_mux u_35_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_36),
    .d1(q_34_37),
    .q(q_35_37)
  );
  

  flop_with_mux u_35_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_37),
    .d1(q_34_38),
    .q(q_35_38)
  );
  

  flop_with_mux u_35_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_35_38),
    .d1(q_34_39),
    .q(q_35_39)
  );
  

  flop_with_mux u_36_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_minus1),
    .d1(q_35_0),
    .q(q_36_0)
  );
  

  flop_with_mux u_36_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_0),
    .d1(q_35_1),
    .q(q_36_1)
  );
  

  flop_with_mux u_36_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_1),
    .d1(q_35_2),
    .q(q_36_2)
  );
  

  flop_with_mux u_36_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_2),
    .d1(q_35_3),
    .q(q_36_3)
  );
  

  flop_with_mux u_36_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_3),
    .d1(q_35_4),
    .q(q_36_4)
  );
  

  flop_with_mux u_36_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_4),
    .d1(q_35_5),
    .q(q_36_5)
  );
  

  flop_with_mux u_36_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_5),
    .d1(q_35_6),
    .q(q_36_6)
  );
  

  flop_with_mux u_36_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_6),
    .d1(q_35_7),
    .q(q_36_7)
  );
  

  flop_with_mux u_36_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_7),
    .d1(q_35_8),
    .q(q_36_8)
  );
  

  flop_with_mux u_36_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_8),
    .d1(q_35_9),
    .q(q_36_9)
  );
  

  flop_with_mux u_36_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_9),
    .d1(q_35_10),
    .q(q_36_10)
  );
  

  flop_with_mux u_36_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_10),
    .d1(q_35_11),
    .q(q_36_11)
  );
  

  flop_with_mux u_36_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_11),
    .d1(q_35_12),
    .q(q_36_12)
  );
  

  flop_with_mux u_36_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_12),
    .d1(q_35_13),
    .q(q_36_13)
  );
  

  flop_with_mux u_36_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_13),
    .d1(q_35_14),
    .q(q_36_14)
  );
  

  flop_with_mux u_36_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_14),
    .d1(q_35_15),
    .q(q_36_15)
  );
  

  flop_with_mux u_36_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_15),
    .d1(q_35_16),
    .q(q_36_16)
  );
  

  flop_with_mux u_36_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_16),
    .d1(q_35_17),
    .q(q_36_17)
  );
  

  flop_with_mux u_36_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_17),
    .d1(q_35_18),
    .q(q_36_18)
  );
  

  flop_with_mux u_36_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_18),
    .d1(q_35_19),
    .q(q_36_19)
  );
  

  flop_with_mux u_36_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_19),
    .d1(q_35_20),
    .q(q_36_20)
  );
  

  flop_with_mux u_36_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_20),
    .d1(q_35_21),
    .q(q_36_21)
  );
  

  flop_with_mux u_36_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_21),
    .d1(q_35_22),
    .q(q_36_22)
  );
  

  flop_with_mux u_36_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_22),
    .d1(q_35_23),
    .q(q_36_23)
  );
  

  flop_with_mux u_36_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_23),
    .d1(q_35_24),
    .q(q_36_24)
  );
  

  flop_with_mux u_36_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_24),
    .d1(q_35_25),
    .q(q_36_25)
  );
  

  flop_with_mux u_36_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_25),
    .d1(q_35_26),
    .q(q_36_26)
  );
  

  flop_with_mux u_36_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_26),
    .d1(q_35_27),
    .q(q_36_27)
  );
  

  flop_with_mux u_36_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_27),
    .d1(q_35_28),
    .q(q_36_28)
  );
  

  flop_with_mux u_36_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_28),
    .d1(q_35_29),
    .q(q_36_29)
  );
  

  flop_with_mux u_36_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_29),
    .d1(q_35_30),
    .q(q_36_30)
  );
  

  flop_with_mux u_36_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_30),
    .d1(q_35_31),
    .q(q_36_31)
  );
  

  flop_with_mux u_36_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_31),
    .d1(q_35_32),
    .q(q_36_32)
  );
  

  flop_with_mux u_36_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_32),
    .d1(q_35_33),
    .q(q_36_33)
  );
  

  flop_with_mux u_36_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_33),
    .d1(q_35_34),
    .q(q_36_34)
  );
  

  flop_with_mux u_36_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_34),
    .d1(q_35_35),
    .q(q_36_35)
  );
  

  flop_with_mux u_36_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_35),
    .d1(q_35_36),
    .q(q_36_36)
  );
  

  flop_with_mux u_36_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_36),
    .d1(q_35_37),
    .q(q_36_37)
  );
  

  flop_with_mux u_36_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_37),
    .d1(q_35_38),
    .q(q_36_38)
  );
  

  flop_with_mux u_36_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_36_38),
    .d1(q_35_39),
    .q(q_36_39)
  );
  

  flop_with_mux u_37_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_minus1),
    .d1(q_36_0),
    .q(q_37_0)
  );
  

  flop_with_mux u_37_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_0),
    .d1(q_36_1),
    .q(q_37_1)
  );
  

  flop_with_mux u_37_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_1),
    .d1(q_36_2),
    .q(q_37_2)
  );
  

  flop_with_mux u_37_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_2),
    .d1(q_36_3),
    .q(q_37_3)
  );
  

  flop_with_mux u_37_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_3),
    .d1(q_36_4),
    .q(q_37_4)
  );
  

  flop_with_mux u_37_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_4),
    .d1(q_36_5),
    .q(q_37_5)
  );
  

  flop_with_mux u_37_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_5),
    .d1(q_36_6),
    .q(q_37_6)
  );
  

  flop_with_mux u_37_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_6),
    .d1(q_36_7),
    .q(q_37_7)
  );
  

  flop_with_mux u_37_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_7),
    .d1(q_36_8),
    .q(q_37_8)
  );
  

  flop_with_mux u_37_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_8),
    .d1(q_36_9),
    .q(q_37_9)
  );
  

  flop_with_mux u_37_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_9),
    .d1(q_36_10),
    .q(q_37_10)
  );
  

  flop_with_mux u_37_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_10),
    .d1(q_36_11),
    .q(q_37_11)
  );
  

  flop_with_mux u_37_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_11),
    .d1(q_36_12),
    .q(q_37_12)
  );
  

  flop_with_mux u_37_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_12),
    .d1(q_36_13),
    .q(q_37_13)
  );
  

  flop_with_mux u_37_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_13),
    .d1(q_36_14),
    .q(q_37_14)
  );
  

  flop_with_mux u_37_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_14),
    .d1(q_36_15),
    .q(q_37_15)
  );
  

  flop_with_mux u_37_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_15),
    .d1(q_36_16),
    .q(q_37_16)
  );
  

  flop_with_mux u_37_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_16),
    .d1(q_36_17),
    .q(q_37_17)
  );
  

  flop_with_mux u_37_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_17),
    .d1(q_36_18),
    .q(q_37_18)
  );
  

  flop_with_mux u_37_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_18),
    .d1(q_36_19),
    .q(q_37_19)
  );
  

  flop_with_mux u_37_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_19),
    .d1(q_36_20),
    .q(q_37_20)
  );
  

  flop_with_mux u_37_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_20),
    .d1(q_36_21),
    .q(q_37_21)
  );
  

  flop_with_mux u_37_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_21),
    .d1(q_36_22),
    .q(q_37_22)
  );
  

  flop_with_mux u_37_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_22),
    .d1(q_36_23),
    .q(q_37_23)
  );
  

  flop_with_mux u_37_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_23),
    .d1(q_36_24),
    .q(q_37_24)
  );
  

  flop_with_mux u_37_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_24),
    .d1(q_36_25),
    .q(q_37_25)
  );
  

  flop_with_mux u_37_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_25),
    .d1(q_36_26),
    .q(q_37_26)
  );
  

  flop_with_mux u_37_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_26),
    .d1(q_36_27),
    .q(q_37_27)
  );
  

  flop_with_mux u_37_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_27),
    .d1(q_36_28),
    .q(q_37_28)
  );
  

  flop_with_mux u_37_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_28),
    .d1(q_36_29),
    .q(q_37_29)
  );
  

  flop_with_mux u_37_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_29),
    .d1(q_36_30),
    .q(q_37_30)
  );
  

  flop_with_mux u_37_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_30),
    .d1(q_36_31),
    .q(q_37_31)
  );
  

  flop_with_mux u_37_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_31),
    .d1(q_36_32),
    .q(q_37_32)
  );
  

  flop_with_mux u_37_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_32),
    .d1(q_36_33),
    .q(q_37_33)
  );
  

  flop_with_mux u_37_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_33),
    .d1(q_36_34),
    .q(q_37_34)
  );
  

  flop_with_mux u_37_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_34),
    .d1(q_36_35),
    .q(q_37_35)
  );
  

  flop_with_mux u_37_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_35),
    .d1(q_36_36),
    .q(q_37_36)
  );
  

  flop_with_mux u_37_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_36),
    .d1(q_36_37),
    .q(q_37_37)
  );
  

  flop_with_mux u_37_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_37),
    .d1(q_36_38),
    .q(q_37_38)
  );
  

  flop_with_mux u_37_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_37_38),
    .d1(q_36_39),
    .q(q_37_39)
  );
  

  flop_with_mux u_38_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_minus1),
    .d1(q_37_0),
    .q(q_38_0)
  );
  

  flop_with_mux u_38_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_0),
    .d1(q_37_1),
    .q(q_38_1)
  );
  

  flop_with_mux u_38_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_1),
    .d1(q_37_2),
    .q(q_38_2)
  );
  

  flop_with_mux u_38_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_2),
    .d1(q_37_3),
    .q(q_38_3)
  );
  

  flop_with_mux u_38_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_3),
    .d1(q_37_4),
    .q(q_38_4)
  );
  

  flop_with_mux u_38_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_4),
    .d1(q_37_5),
    .q(q_38_5)
  );
  

  flop_with_mux u_38_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_5),
    .d1(q_37_6),
    .q(q_38_6)
  );
  

  flop_with_mux u_38_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_6),
    .d1(q_37_7),
    .q(q_38_7)
  );
  

  flop_with_mux u_38_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_7),
    .d1(q_37_8),
    .q(q_38_8)
  );
  

  flop_with_mux u_38_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_8),
    .d1(q_37_9),
    .q(q_38_9)
  );
  

  flop_with_mux u_38_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_9),
    .d1(q_37_10),
    .q(q_38_10)
  );
  

  flop_with_mux u_38_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_10),
    .d1(q_37_11),
    .q(q_38_11)
  );
  

  flop_with_mux u_38_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_11),
    .d1(q_37_12),
    .q(q_38_12)
  );
  

  flop_with_mux u_38_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_12),
    .d1(q_37_13),
    .q(q_38_13)
  );
  

  flop_with_mux u_38_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_13),
    .d1(q_37_14),
    .q(q_38_14)
  );
  

  flop_with_mux u_38_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_14),
    .d1(q_37_15),
    .q(q_38_15)
  );
  

  flop_with_mux u_38_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_15),
    .d1(q_37_16),
    .q(q_38_16)
  );
  

  flop_with_mux u_38_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_16),
    .d1(q_37_17),
    .q(q_38_17)
  );
  

  flop_with_mux u_38_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_17),
    .d1(q_37_18),
    .q(q_38_18)
  );
  

  flop_with_mux u_38_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_18),
    .d1(q_37_19),
    .q(q_38_19)
  );
  

  flop_with_mux u_38_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_19),
    .d1(q_37_20),
    .q(q_38_20)
  );
  

  flop_with_mux u_38_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_20),
    .d1(q_37_21),
    .q(q_38_21)
  );
  

  flop_with_mux u_38_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_21),
    .d1(q_37_22),
    .q(q_38_22)
  );
  

  flop_with_mux u_38_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_22),
    .d1(q_37_23),
    .q(q_38_23)
  );
  

  flop_with_mux u_38_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_23),
    .d1(q_37_24),
    .q(q_38_24)
  );
  

  flop_with_mux u_38_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_24),
    .d1(q_37_25),
    .q(q_38_25)
  );
  

  flop_with_mux u_38_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_25),
    .d1(q_37_26),
    .q(q_38_26)
  );
  

  flop_with_mux u_38_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_26),
    .d1(q_37_27),
    .q(q_38_27)
  );
  

  flop_with_mux u_38_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_27),
    .d1(q_37_28),
    .q(q_38_28)
  );
  

  flop_with_mux u_38_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_28),
    .d1(q_37_29),
    .q(q_38_29)
  );
  

  flop_with_mux u_38_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_29),
    .d1(q_37_30),
    .q(q_38_30)
  );
  

  flop_with_mux u_38_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_30),
    .d1(q_37_31),
    .q(q_38_31)
  );
  

  flop_with_mux u_38_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_31),
    .d1(q_37_32),
    .q(q_38_32)
  );
  

  flop_with_mux u_38_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_32),
    .d1(q_37_33),
    .q(q_38_33)
  );
  

  flop_with_mux u_38_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_33),
    .d1(q_37_34),
    .q(q_38_34)
  );
  

  flop_with_mux u_38_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_34),
    .d1(q_37_35),
    .q(q_38_35)
  );
  

  flop_with_mux u_38_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_35),
    .d1(q_37_36),
    .q(q_38_36)
  );
  

  flop_with_mux u_38_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_36),
    .d1(q_37_37),
    .q(q_38_37)
  );
  

  flop_with_mux u_38_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_37),
    .d1(q_37_38),
    .q(q_38_38)
  );
  

  flop_with_mux u_38_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_38_38),
    .d1(q_37_39),
    .q(q_38_39)
  );
  

  flop_with_mux u_39_0 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_minus1),
    .d1(q_38_0),
    .q(q_39_0)
  );
  

  flop_with_mux u_39_1 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_0),
    .d1(q_38_1),
    .q(q_39_1)
  );
  

  flop_with_mux u_39_2 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_1),
    .d1(q_38_2),
    .q(q_39_2)
  );
  

  flop_with_mux u_39_3 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_2),
    .d1(q_38_3),
    .q(q_39_3)
  );
  

  flop_with_mux u_39_4 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_3),
    .d1(q_38_4),
    .q(q_39_4)
  );
  

  flop_with_mux u_39_5 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_4),
    .d1(q_38_5),
    .q(q_39_5)
  );
  

  flop_with_mux u_39_6 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_5),
    .d1(q_38_6),
    .q(q_39_6)
  );
  

  flop_with_mux u_39_7 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_6),
    .d1(q_38_7),
    .q(q_39_7)
  );
  

  flop_with_mux u_39_8 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_7),
    .d1(q_38_8),
    .q(q_39_8)
  );
  

  flop_with_mux u_39_9 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_8),
    .d1(q_38_9),
    .q(q_39_9)
  );
  

  flop_with_mux u_39_10 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_9),
    .d1(q_38_10),
    .q(q_39_10)
  );
  

  flop_with_mux u_39_11 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_10),
    .d1(q_38_11),
    .q(q_39_11)
  );
  

  flop_with_mux u_39_12 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_11),
    .d1(q_38_12),
    .q(q_39_12)
  );
  

  flop_with_mux u_39_13 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_12),
    .d1(q_38_13),
    .q(q_39_13)
  );
  

  flop_with_mux u_39_14 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_13),
    .d1(q_38_14),
    .q(q_39_14)
  );
  

  flop_with_mux u_39_15 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_14),
    .d1(q_38_15),
    .q(q_39_15)
  );
  

  flop_with_mux u_39_16 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_15),
    .d1(q_38_16),
    .q(q_39_16)
  );
  

  flop_with_mux u_39_17 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_16),
    .d1(q_38_17),
    .q(q_39_17)
  );
  

  flop_with_mux u_39_18 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_17),
    .d1(q_38_18),
    .q(q_39_18)
  );
  

  flop_with_mux u_39_19 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_18),
    .d1(q_38_19),
    .q(q_39_19)
  );
  

  flop_with_mux u_39_20 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_19),
    .d1(q_38_20),
    .q(q_39_20)
  );
  

  flop_with_mux u_39_21 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_20),
    .d1(q_38_21),
    .q(q_39_21)
  );
  

  flop_with_mux u_39_22 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_21),
    .d1(q_38_22),
    .q(q_39_22)
  );
  

  flop_with_mux u_39_23 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_22),
    .d1(q_38_23),
    .q(q_39_23)
  );
  

  flop_with_mux u_39_24 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_23),
    .d1(q_38_24),
    .q(q_39_24)
  );
  

  flop_with_mux u_39_25 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_24),
    .d1(q_38_25),
    .q(q_39_25)
  );
  

  flop_with_mux u_39_26 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_25),
    .d1(q_38_26),
    .q(q_39_26)
  );
  

  flop_with_mux u_39_27 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_26),
    .d1(q_38_27),
    .q(q_39_27)
  );
  

  flop_with_mux u_39_28 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_27),
    .d1(q_38_28),
    .q(q_39_28)
  );
  

  flop_with_mux u_39_29 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_28),
    .d1(q_38_29),
    .q(q_39_29)
  );
  

  flop_with_mux u_39_30 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_29),
    .d1(q_38_30),
    .q(q_39_30)
  );
  

  flop_with_mux u_39_31 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_30),
    .d1(q_38_31),
    .q(q_39_31)
  );
  

  flop_with_mux u_39_32 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_31),
    .d1(q_38_32),
    .q(q_39_32)
  );
  

  flop_with_mux u_39_33 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_32),
    .d1(q_38_33),
    .q(q_39_33)
  );
  

  flop_with_mux u_39_34 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_33),
    .d1(q_38_34),
    .q(q_39_34)
  );
  

  flop_with_mux u_39_35 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_34),
    .d1(q_38_35),
    .q(q_39_35)
  );
  

  flop_with_mux u_39_36 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_35),
    .d1(q_38_36),
    .q(q_39_36)
  );
  

  flop_with_mux u_39_37 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_36),
    .d1(q_38_37),
    .q(q_39_37)
  );
  

  flop_with_mux u_39_38 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_37),
    .d1(q_38_38),
    .q(q_39_38)
  );
  

  flop_with_mux u_39_39 (
    .clk(clk),
    .valid(valid),
    .sel(load_unload), //0 for load (left to right), 1 for unload (top to bottom)
    .d0(q_39_38),
    .d1(q_38_39),
    .q(q_39_39)
  );
  
endmodule

